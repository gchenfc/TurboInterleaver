
library ieee;
use ieee.std_logic_1164.all;

entity TurboInterleaver_Interleaver is
	port (
		clk, reset_async:			in std_logic;

		dataBufferIn_short:			in std_logic_vector(1055 DOWNTO 0);
		dataBufferIn_long:			in std_logic_vector(6143 DOWNTO 0);
		dataBufferOut_short:		out std_logic_vector(1055 DOWNTO 0);
		dataBufferOut_long:			out std_logic_vector(6143 DOWNTO 0)
	);
end TurboInterleaver_Interleaver;

architecture arch1 of TurboInterleaver_Interleaver is

begin

	dataBufferOut_short(   0) <= dataBufferIn_short(   0);
	dataBufferOut_short(  83) <= dataBufferIn_short(   1);
	dataBufferOut_short( 166) <= dataBufferIn_short(   2);
	dataBufferOut_short( 249) <= dataBufferIn_short(   3);
	dataBufferOut_short( 332) <= dataBufferIn_short(   4);
	dataBufferOut_short( 415) <= dataBufferIn_short(   5);
	dataBufferOut_short( 498) <= dataBufferIn_short(   6);
	dataBufferOut_short( 581) <= dataBufferIn_short(   7);
	dataBufferOut_short( 664) <= dataBufferIn_short(   8);
	dataBufferOut_short( 747) <= dataBufferIn_short(   9);
	dataBufferOut_short( 830) <= dataBufferIn_short(  10);
	dataBufferOut_short( 913) <= dataBufferIn_short(  11);
	dataBufferOut_short( 996) <= dataBufferIn_short(  12);
	dataBufferOut_short(  23) <= dataBufferIn_short(  13);
	dataBufferOut_short( 106) <= dataBufferIn_short(  14);
	dataBufferOut_short( 189) <= dataBufferIn_short(  15);
	dataBufferOut_short( 272) <= dataBufferIn_short(  16);
	dataBufferOut_short( 355) <= dataBufferIn_short(  17);
	dataBufferOut_short( 438) <= dataBufferIn_short(  18);
	dataBufferOut_short( 521) <= dataBufferIn_short(  19);
	dataBufferOut_short( 604) <= dataBufferIn_short(  20);
	dataBufferOut_short( 687) <= dataBufferIn_short(  21);
	dataBufferOut_short( 770) <= dataBufferIn_short(  22);
	dataBufferOut_short( 853) <= dataBufferIn_short(  23);
	dataBufferOut_short( 936) <= dataBufferIn_short(  24);
	dataBufferOut_short(1019) <= dataBufferIn_short(  25);
	dataBufferOut_short(  46) <= dataBufferIn_short(  26);
	dataBufferOut_short( 129) <= dataBufferIn_short(  27);
	dataBufferOut_short( 212) <= dataBufferIn_short(  28);
	dataBufferOut_short( 295) <= dataBufferIn_short(  29);
	dataBufferOut_short( 378) <= dataBufferIn_short(  30);
	dataBufferOut_short( 461) <= dataBufferIn_short(  31);
	dataBufferOut_short( 544) <= dataBufferIn_short(  32);
	dataBufferOut_short( 627) <= dataBufferIn_short(  33);
	dataBufferOut_short( 710) <= dataBufferIn_short(  34);
	dataBufferOut_short( 793) <= dataBufferIn_short(  35);
	dataBufferOut_short( 876) <= dataBufferIn_short(  36);
	dataBufferOut_short( 959) <= dataBufferIn_short(  37);
	dataBufferOut_short(1042) <= dataBufferIn_short(  38);
	dataBufferOut_short(  69) <= dataBufferIn_short(  39);
	dataBufferOut_short( 152) <= dataBufferIn_short(  40);
	dataBufferOut_short( 235) <= dataBufferIn_short(  41);
	dataBufferOut_short( 318) <= dataBufferIn_short(  42);
	dataBufferOut_short( 401) <= dataBufferIn_short(  43);
	dataBufferOut_short( 484) <= dataBufferIn_short(  44);
	dataBufferOut_short( 567) <= dataBufferIn_short(  45);
	dataBufferOut_short( 650) <= dataBufferIn_short(  46);
	dataBufferOut_short( 733) <= dataBufferIn_short(  47);
	dataBufferOut_short( 816) <= dataBufferIn_short(  48);
	dataBufferOut_short( 899) <= dataBufferIn_short(  49);
	dataBufferOut_short( 982) <= dataBufferIn_short(  50);
	dataBufferOut_short(   9) <= dataBufferIn_short(  51);
	dataBufferOut_short(  92) <= dataBufferIn_short(  52);
	dataBufferOut_short( 175) <= dataBufferIn_short(  53);
	dataBufferOut_short( 258) <= dataBufferIn_short(  54);
	dataBufferOut_short( 341) <= dataBufferIn_short(  55);
	dataBufferOut_short( 424) <= dataBufferIn_short(  56);
	dataBufferOut_short( 507) <= dataBufferIn_short(  57);
	dataBufferOut_short( 590) <= dataBufferIn_short(  58);
	dataBufferOut_short( 673) <= dataBufferIn_short(  59);
	dataBufferOut_short( 756) <= dataBufferIn_short(  60);
	dataBufferOut_short( 839) <= dataBufferIn_short(  61);
	dataBufferOut_short( 922) <= dataBufferIn_short(  62);
	dataBufferOut_short(1005) <= dataBufferIn_short(  63);
	dataBufferOut_short(  32) <= dataBufferIn_short(  64);
	dataBufferOut_short( 115) <= dataBufferIn_short(  65);
	dataBufferOut_short( 198) <= dataBufferIn_short(  66);
	dataBufferOut_short( 281) <= dataBufferIn_short(  67);
	dataBufferOut_short( 364) <= dataBufferIn_short(  68);
	dataBufferOut_short( 447) <= dataBufferIn_short(  69);
	dataBufferOut_short( 530) <= dataBufferIn_short(  70);
	dataBufferOut_short( 613) <= dataBufferIn_short(  71);
	dataBufferOut_short( 696) <= dataBufferIn_short(  72);
	dataBufferOut_short( 779) <= dataBufferIn_short(  73);
	dataBufferOut_short( 862) <= dataBufferIn_short(  74);
	dataBufferOut_short( 945) <= dataBufferIn_short(  75);
	dataBufferOut_short(1028) <= dataBufferIn_short(  76);
	dataBufferOut_short(  55) <= dataBufferIn_short(  77);
	dataBufferOut_short( 138) <= dataBufferIn_short(  78);
	dataBufferOut_short( 221) <= dataBufferIn_short(  79);
	dataBufferOut_short( 304) <= dataBufferIn_short(  80);
	dataBufferOut_short( 387) <= dataBufferIn_short(  81);
	dataBufferOut_short( 470) <= dataBufferIn_short(  82);
	dataBufferOut_short( 553) <= dataBufferIn_short(  83);
	dataBufferOut_short( 636) <= dataBufferIn_short(  84);
	dataBufferOut_short( 719) <= dataBufferIn_short(  85);
	dataBufferOut_short( 802) <= dataBufferIn_short(  86);
	dataBufferOut_short( 885) <= dataBufferIn_short(  87);
	dataBufferOut_short( 968) <= dataBufferIn_short(  88);
	dataBufferOut_short(1051) <= dataBufferIn_short(  89);
	dataBufferOut_short(  78) <= dataBufferIn_short(  90);
	dataBufferOut_short( 161) <= dataBufferIn_short(  91);
	dataBufferOut_short( 244) <= dataBufferIn_short(  92);
	dataBufferOut_short( 327) <= dataBufferIn_short(  93);
	dataBufferOut_short( 410) <= dataBufferIn_short(  94);
	dataBufferOut_short( 493) <= dataBufferIn_short(  95);
	dataBufferOut_short( 576) <= dataBufferIn_short(  96);
	dataBufferOut_short( 659) <= dataBufferIn_short(  97);
	dataBufferOut_short( 742) <= dataBufferIn_short(  98);
	dataBufferOut_short( 825) <= dataBufferIn_short(  99);
	dataBufferOut_short( 908) <= dataBufferIn_short( 100);
	dataBufferOut_short( 991) <= dataBufferIn_short( 101);
	dataBufferOut_short(  18) <= dataBufferIn_short( 102);
	dataBufferOut_short( 101) <= dataBufferIn_short( 103);
	dataBufferOut_short( 184) <= dataBufferIn_short( 104);
	dataBufferOut_short( 267) <= dataBufferIn_short( 105);
	dataBufferOut_short( 350) <= dataBufferIn_short( 106);
	dataBufferOut_short( 433) <= dataBufferIn_short( 107);
	dataBufferOut_short( 516) <= dataBufferIn_short( 108);
	dataBufferOut_short( 599) <= dataBufferIn_short( 109);
	dataBufferOut_short( 682) <= dataBufferIn_short( 110);
	dataBufferOut_short( 765) <= dataBufferIn_short( 111);
	dataBufferOut_short( 848) <= dataBufferIn_short( 112);
	dataBufferOut_short( 931) <= dataBufferIn_short( 113);
	dataBufferOut_short(1014) <= dataBufferIn_short( 114);
	dataBufferOut_short(  41) <= dataBufferIn_short( 115);
	dataBufferOut_short( 124) <= dataBufferIn_short( 116);
	dataBufferOut_short( 207) <= dataBufferIn_short( 117);
	dataBufferOut_short( 290) <= dataBufferIn_short( 118);
	dataBufferOut_short( 373) <= dataBufferIn_short( 119);
	dataBufferOut_short( 456) <= dataBufferIn_short( 120);
	dataBufferOut_short( 539) <= dataBufferIn_short( 121);
	dataBufferOut_short( 622) <= dataBufferIn_short( 122);
	dataBufferOut_short( 705) <= dataBufferIn_short( 123);
	dataBufferOut_short( 788) <= dataBufferIn_short( 124);
	dataBufferOut_short( 871) <= dataBufferIn_short( 125);
	dataBufferOut_short( 954) <= dataBufferIn_short( 126);
	dataBufferOut_short(1037) <= dataBufferIn_short( 127);
	dataBufferOut_short(  64) <= dataBufferIn_short( 128);
	dataBufferOut_short( 147) <= dataBufferIn_short( 129);
	dataBufferOut_short( 230) <= dataBufferIn_short( 130);
	dataBufferOut_short( 313) <= dataBufferIn_short( 131);
	dataBufferOut_short( 396) <= dataBufferIn_short( 132);
	dataBufferOut_short( 479) <= dataBufferIn_short( 133);
	dataBufferOut_short( 562) <= dataBufferIn_short( 134);
	dataBufferOut_short( 645) <= dataBufferIn_short( 135);
	dataBufferOut_short( 728) <= dataBufferIn_short( 136);
	dataBufferOut_short( 811) <= dataBufferIn_short( 137);
	dataBufferOut_short( 894) <= dataBufferIn_short( 138);
	dataBufferOut_short( 977) <= dataBufferIn_short( 139);
	dataBufferOut_short(   4) <= dataBufferIn_short( 140);
	dataBufferOut_short(  87) <= dataBufferIn_short( 141);
	dataBufferOut_short( 170) <= dataBufferIn_short( 142);
	dataBufferOut_short( 253) <= dataBufferIn_short( 143);
	dataBufferOut_short( 336) <= dataBufferIn_short( 144);
	dataBufferOut_short( 419) <= dataBufferIn_short( 145);
	dataBufferOut_short( 502) <= dataBufferIn_short( 146);
	dataBufferOut_short( 585) <= dataBufferIn_short( 147);
	dataBufferOut_short( 668) <= dataBufferIn_short( 148);
	dataBufferOut_short( 751) <= dataBufferIn_short( 149);
	dataBufferOut_short( 834) <= dataBufferIn_short( 150);
	dataBufferOut_short( 917) <= dataBufferIn_short( 151);
	dataBufferOut_short(1000) <= dataBufferIn_short( 152);
	dataBufferOut_short(  27) <= dataBufferIn_short( 153);
	dataBufferOut_short( 110) <= dataBufferIn_short( 154);
	dataBufferOut_short( 193) <= dataBufferIn_short( 155);
	dataBufferOut_short( 276) <= dataBufferIn_short( 156);
	dataBufferOut_short( 359) <= dataBufferIn_short( 157);
	dataBufferOut_short( 442) <= dataBufferIn_short( 158);
	dataBufferOut_short( 525) <= dataBufferIn_short( 159);
	dataBufferOut_short( 608) <= dataBufferIn_short( 160);
	dataBufferOut_short( 691) <= dataBufferIn_short( 161);
	dataBufferOut_short( 774) <= dataBufferIn_short( 162);
	dataBufferOut_short( 857) <= dataBufferIn_short( 163);
	dataBufferOut_short( 940) <= dataBufferIn_short( 164);
	dataBufferOut_short(1023) <= dataBufferIn_short( 165);
	dataBufferOut_short(  50) <= dataBufferIn_short( 166);
	dataBufferOut_short( 133) <= dataBufferIn_short( 167);
	dataBufferOut_short( 216) <= dataBufferIn_short( 168);
	dataBufferOut_short( 299) <= dataBufferIn_short( 169);
	dataBufferOut_short( 382) <= dataBufferIn_short( 170);
	dataBufferOut_short( 465) <= dataBufferIn_short( 171);
	dataBufferOut_short( 548) <= dataBufferIn_short( 172);
	dataBufferOut_short( 631) <= dataBufferIn_short( 173);
	dataBufferOut_short( 714) <= dataBufferIn_short( 174);
	dataBufferOut_short( 797) <= dataBufferIn_short( 175);
	dataBufferOut_short( 880) <= dataBufferIn_short( 176);
	dataBufferOut_short( 963) <= dataBufferIn_short( 177);
	dataBufferOut_short(1046) <= dataBufferIn_short( 178);
	dataBufferOut_short(  73) <= dataBufferIn_short( 179);
	dataBufferOut_short( 156) <= dataBufferIn_short( 180);
	dataBufferOut_short( 239) <= dataBufferIn_short( 181);
	dataBufferOut_short( 322) <= dataBufferIn_short( 182);
	dataBufferOut_short( 405) <= dataBufferIn_short( 183);
	dataBufferOut_short( 488) <= dataBufferIn_short( 184);
	dataBufferOut_short( 571) <= dataBufferIn_short( 185);
	dataBufferOut_short( 654) <= dataBufferIn_short( 186);
	dataBufferOut_short( 737) <= dataBufferIn_short( 187);
	dataBufferOut_short( 820) <= dataBufferIn_short( 188);
	dataBufferOut_short( 903) <= dataBufferIn_short( 189);
	dataBufferOut_short( 986) <= dataBufferIn_short( 190);
	dataBufferOut_short(  13) <= dataBufferIn_short( 191);
	dataBufferOut_short(  96) <= dataBufferIn_short( 192);
	dataBufferOut_short( 179) <= dataBufferIn_short( 193);
	dataBufferOut_short( 262) <= dataBufferIn_short( 194);
	dataBufferOut_short( 345) <= dataBufferIn_short( 195);
	dataBufferOut_short( 428) <= dataBufferIn_short( 196);
	dataBufferOut_short( 511) <= dataBufferIn_short( 197);
	dataBufferOut_short( 594) <= dataBufferIn_short( 198);
	dataBufferOut_short( 677) <= dataBufferIn_short( 199);
	dataBufferOut_short( 760) <= dataBufferIn_short( 200);
	dataBufferOut_short( 843) <= dataBufferIn_short( 201);
	dataBufferOut_short( 926) <= dataBufferIn_short( 202);
	dataBufferOut_short(1009) <= dataBufferIn_short( 203);
	dataBufferOut_short(  36) <= dataBufferIn_short( 204);
	dataBufferOut_short( 119) <= dataBufferIn_short( 205);
	dataBufferOut_short( 202) <= dataBufferIn_short( 206);
	dataBufferOut_short( 285) <= dataBufferIn_short( 207);
	dataBufferOut_short( 368) <= dataBufferIn_short( 208);
	dataBufferOut_short( 451) <= dataBufferIn_short( 209);
	dataBufferOut_short( 534) <= dataBufferIn_short( 210);
	dataBufferOut_short( 617) <= dataBufferIn_short( 211);
	dataBufferOut_short( 700) <= dataBufferIn_short( 212);
	dataBufferOut_short( 783) <= dataBufferIn_short( 213);
	dataBufferOut_short( 866) <= dataBufferIn_short( 214);
	dataBufferOut_short( 949) <= dataBufferIn_short( 215);
	dataBufferOut_short(1032) <= dataBufferIn_short( 216);
	dataBufferOut_short(  59) <= dataBufferIn_short( 217);
	dataBufferOut_short( 142) <= dataBufferIn_short( 218);
	dataBufferOut_short( 225) <= dataBufferIn_short( 219);
	dataBufferOut_short( 308) <= dataBufferIn_short( 220);
	dataBufferOut_short( 391) <= dataBufferIn_short( 221);
	dataBufferOut_short( 474) <= dataBufferIn_short( 222);
	dataBufferOut_short( 557) <= dataBufferIn_short( 223);
	dataBufferOut_short( 640) <= dataBufferIn_short( 224);
	dataBufferOut_short( 723) <= dataBufferIn_short( 225);
	dataBufferOut_short( 806) <= dataBufferIn_short( 226);
	dataBufferOut_short( 889) <= dataBufferIn_short( 227);
	dataBufferOut_short( 972) <= dataBufferIn_short( 228);
	dataBufferOut_short(1055) <= dataBufferIn_short( 229);
	dataBufferOut_short(  82) <= dataBufferIn_short( 230);
	dataBufferOut_short( 165) <= dataBufferIn_short( 231);
	dataBufferOut_short( 248) <= dataBufferIn_short( 232);
	dataBufferOut_short( 331) <= dataBufferIn_short( 233);
	dataBufferOut_short( 414) <= dataBufferIn_short( 234);
	dataBufferOut_short( 497) <= dataBufferIn_short( 235);
	dataBufferOut_short( 580) <= dataBufferIn_short( 236);
	dataBufferOut_short( 663) <= dataBufferIn_short( 237);
	dataBufferOut_short( 746) <= dataBufferIn_short( 238);
	dataBufferOut_short( 829) <= dataBufferIn_short( 239);
	dataBufferOut_short( 912) <= dataBufferIn_short( 240);
	dataBufferOut_short( 995) <= dataBufferIn_short( 241);
	dataBufferOut_short(  22) <= dataBufferIn_short( 242);
	dataBufferOut_short( 105) <= dataBufferIn_short( 243);
	dataBufferOut_short( 188) <= dataBufferIn_short( 244);
	dataBufferOut_short( 271) <= dataBufferIn_short( 245);
	dataBufferOut_short( 354) <= dataBufferIn_short( 246);
	dataBufferOut_short( 437) <= dataBufferIn_short( 247);
	dataBufferOut_short( 520) <= dataBufferIn_short( 248);
	dataBufferOut_short( 603) <= dataBufferIn_short( 249);
	dataBufferOut_short( 686) <= dataBufferIn_short( 250);
	dataBufferOut_short( 769) <= dataBufferIn_short( 251);
	dataBufferOut_short( 852) <= dataBufferIn_short( 252);
	dataBufferOut_short( 935) <= dataBufferIn_short( 253);
	dataBufferOut_short(1018) <= dataBufferIn_short( 254);
	dataBufferOut_short(  45) <= dataBufferIn_short( 255);
	dataBufferOut_short( 128) <= dataBufferIn_short( 256);
	dataBufferOut_short( 211) <= dataBufferIn_short( 257);
	dataBufferOut_short( 294) <= dataBufferIn_short( 258);
	dataBufferOut_short( 377) <= dataBufferIn_short( 259);
	dataBufferOut_short( 460) <= dataBufferIn_short( 260);
	dataBufferOut_short( 543) <= dataBufferIn_short( 261);
	dataBufferOut_short( 626) <= dataBufferIn_short( 262);
	dataBufferOut_short( 709) <= dataBufferIn_short( 263);
	dataBufferOut_short( 792) <= dataBufferIn_short( 264);
	dataBufferOut_short( 875) <= dataBufferIn_short( 265);
	dataBufferOut_short( 958) <= dataBufferIn_short( 266);
	dataBufferOut_short(1041) <= dataBufferIn_short( 267);
	dataBufferOut_short(  68) <= dataBufferIn_short( 268);
	dataBufferOut_short( 151) <= dataBufferIn_short( 269);
	dataBufferOut_short( 234) <= dataBufferIn_short( 270);
	dataBufferOut_short( 317) <= dataBufferIn_short( 271);
	dataBufferOut_short( 400) <= dataBufferIn_short( 272);
	dataBufferOut_short( 483) <= dataBufferIn_short( 273);
	dataBufferOut_short( 566) <= dataBufferIn_short( 274);
	dataBufferOut_short( 649) <= dataBufferIn_short( 275);
	dataBufferOut_short( 732) <= dataBufferIn_short( 276);
	dataBufferOut_short( 815) <= dataBufferIn_short( 277);
	dataBufferOut_short( 898) <= dataBufferIn_short( 278);
	dataBufferOut_short( 981) <= dataBufferIn_short( 279);
	dataBufferOut_short(   8) <= dataBufferIn_short( 280);
	dataBufferOut_short(  91) <= dataBufferIn_short( 281);
	dataBufferOut_short( 174) <= dataBufferIn_short( 282);
	dataBufferOut_short( 257) <= dataBufferIn_short( 283);
	dataBufferOut_short( 340) <= dataBufferIn_short( 284);
	dataBufferOut_short( 423) <= dataBufferIn_short( 285);
	dataBufferOut_short( 506) <= dataBufferIn_short( 286);
	dataBufferOut_short( 589) <= dataBufferIn_short( 287);
	dataBufferOut_short( 672) <= dataBufferIn_short( 288);
	dataBufferOut_short( 755) <= dataBufferIn_short( 289);
	dataBufferOut_short( 838) <= dataBufferIn_short( 290);
	dataBufferOut_short( 921) <= dataBufferIn_short( 291);
	dataBufferOut_short(1004) <= dataBufferIn_short( 292);
	dataBufferOut_short(  31) <= dataBufferIn_short( 293);
	dataBufferOut_short( 114) <= dataBufferIn_short( 294);
	dataBufferOut_short( 197) <= dataBufferIn_short( 295);
	dataBufferOut_short( 280) <= dataBufferIn_short( 296);
	dataBufferOut_short( 363) <= dataBufferIn_short( 297);
	dataBufferOut_short( 446) <= dataBufferIn_short( 298);
	dataBufferOut_short( 529) <= dataBufferIn_short( 299);
	dataBufferOut_short( 612) <= dataBufferIn_short( 300);
	dataBufferOut_short( 695) <= dataBufferIn_short( 301);
	dataBufferOut_short( 778) <= dataBufferIn_short( 302);
	dataBufferOut_short( 861) <= dataBufferIn_short( 303);
	dataBufferOut_short( 944) <= dataBufferIn_short( 304);
	dataBufferOut_short(1027) <= dataBufferIn_short( 305);
	dataBufferOut_short(  54) <= dataBufferIn_short( 306);
	dataBufferOut_short( 137) <= dataBufferIn_short( 307);
	dataBufferOut_short( 220) <= dataBufferIn_short( 308);
	dataBufferOut_short( 303) <= dataBufferIn_short( 309);
	dataBufferOut_short( 386) <= dataBufferIn_short( 310);
	dataBufferOut_short( 469) <= dataBufferIn_short( 311);
	dataBufferOut_short( 552) <= dataBufferIn_short( 312);
	dataBufferOut_short( 635) <= dataBufferIn_short( 313);
	dataBufferOut_short( 718) <= dataBufferIn_short( 314);
	dataBufferOut_short( 801) <= dataBufferIn_short( 315);
	dataBufferOut_short( 884) <= dataBufferIn_short( 316);
	dataBufferOut_short( 967) <= dataBufferIn_short( 317);
	dataBufferOut_short(1050) <= dataBufferIn_short( 318);
	dataBufferOut_short(  77) <= dataBufferIn_short( 319);
	dataBufferOut_short( 160) <= dataBufferIn_short( 320);
	dataBufferOut_short( 243) <= dataBufferIn_short( 321);
	dataBufferOut_short( 326) <= dataBufferIn_short( 322);
	dataBufferOut_short( 409) <= dataBufferIn_short( 323);
	dataBufferOut_short( 492) <= dataBufferIn_short( 324);
	dataBufferOut_short( 575) <= dataBufferIn_short( 325);
	dataBufferOut_short( 658) <= dataBufferIn_short( 326);
	dataBufferOut_short( 741) <= dataBufferIn_short( 327);
	dataBufferOut_short( 824) <= dataBufferIn_short( 328);
	dataBufferOut_short( 907) <= dataBufferIn_short( 329);
	dataBufferOut_short( 990) <= dataBufferIn_short( 330);
	dataBufferOut_short(  17) <= dataBufferIn_short( 331);
	dataBufferOut_short( 100) <= dataBufferIn_short( 332);
	dataBufferOut_short( 183) <= dataBufferIn_short( 333);
	dataBufferOut_short( 266) <= dataBufferIn_short( 334);
	dataBufferOut_short( 349) <= dataBufferIn_short( 335);
	dataBufferOut_short( 432) <= dataBufferIn_short( 336);
	dataBufferOut_short( 515) <= dataBufferIn_short( 337);
	dataBufferOut_short( 598) <= dataBufferIn_short( 338);
	dataBufferOut_short( 681) <= dataBufferIn_short( 339);
	dataBufferOut_short( 764) <= dataBufferIn_short( 340);
	dataBufferOut_short( 847) <= dataBufferIn_short( 341);
	dataBufferOut_short( 930) <= dataBufferIn_short( 342);
	dataBufferOut_short(1013) <= dataBufferIn_short( 343);
	dataBufferOut_short(  40) <= dataBufferIn_short( 344);
	dataBufferOut_short( 123) <= dataBufferIn_short( 345);
	dataBufferOut_short( 206) <= dataBufferIn_short( 346);
	dataBufferOut_short( 289) <= dataBufferIn_short( 347);
	dataBufferOut_short( 372) <= dataBufferIn_short( 348);
	dataBufferOut_short( 455) <= dataBufferIn_short( 349);
	dataBufferOut_short( 538) <= dataBufferIn_short( 350);
	dataBufferOut_short( 621) <= dataBufferIn_short( 351);
	dataBufferOut_short( 704) <= dataBufferIn_short( 352);
	dataBufferOut_short( 787) <= dataBufferIn_short( 353);
	dataBufferOut_short( 870) <= dataBufferIn_short( 354);
	dataBufferOut_short( 953) <= dataBufferIn_short( 355);
	dataBufferOut_short(1036) <= dataBufferIn_short( 356);
	dataBufferOut_short(  63) <= dataBufferIn_short( 357);
	dataBufferOut_short( 146) <= dataBufferIn_short( 358);
	dataBufferOut_short( 229) <= dataBufferIn_short( 359);
	dataBufferOut_short( 312) <= dataBufferIn_short( 360);
	dataBufferOut_short( 395) <= dataBufferIn_short( 361);
	dataBufferOut_short( 478) <= dataBufferIn_short( 362);
	dataBufferOut_short( 561) <= dataBufferIn_short( 363);
	dataBufferOut_short( 644) <= dataBufferIn_short( 364);
	dataBufferOut_short( 727) <= dataBufferIn_short( 365);
	dataBufferOut_short( 810) <= dataBufferIn_short( 366);
	dataBufferOut_short( 893) <= dataBufferIn_short( 367);
	dataBufferOut_short( 976) <= dataBufferIn_short( 368);
	dataBufferOut_short(   3) <= dataBufferIn_short( 369);
	dataBufferOut_short(  86) <= dataBufferIn_short( 370);
	dataBufferOut_short( 169) <= dataBufferIn_short( 371);
	dataBufferOut_short( 252) <= dataBufferIn_short( 372);
	dataBufferOut_short( 335) <= dataBufferIn_short( 373);
	dataBufferOut_short( 418) <= dataBufferIn_short( 374);
	dataBufferOut_short( 501) <= dataBufferIn_short( 375);
	dataBufferOut_short( 584) <= dataBufferIn_short( 376);
	dataBufferOut_short( 667) <= dataBufferIn_short( 377);
	dataBufferOut_short( 750) <= dataBufferIn_short( 378);
	dataBufferOut_short( 833) <= dataBufferIn_short( 379);
	dataBufferOut_short( 916) <= dataBufferIn_short( 380);
	dataBufferOut_short( 999) <= dataBufferIn_short( 381);
	dataBufferOut_short(  26) <= dataBufferIn_short( 382);
	dataBufferOut_short( 109) <= dataBufferIn_short( 383);
	dataBufferOut_short( 192) <= dataBufferIn_short( 384);
	dataBufferOut_short( 275) <= dataBufferIn_short( 385);
	dataBufferOut_short( 358) <= dataBufferIn_short( 386);
	dataBufferOut_short( 441) <= dataBufferIn_short( 387);
	dataBufferOut_short( 524) <= dataBufferIn_short( 388);
	dataBufferOut_short( 607) <= dataBufferIn_short( 389);
	dataBufferOut_short( 690) <= dataBufferIn_short( 390);
	dataBufferOut_short( 773) <= dataBufferIn_short( 391);
	dataBufferOut_short( 856) <= dataBufferIn_short( 392);
	dataBufferOut_short( 939) <= dataBufferIn_short( 393);
	dataBufferOut_short(1022) <= dataBufferIn_short( 394);
	dataBufferOut_short(  49) <= dataBufferIn_short( 395);
	dataBufferOut_short( 132) <= dataBufferIn_short( 396);
	dataBufferOut_short( 215) <= dataBufferIn_short( 397);
	dataBufferOut_short( 298) <= dataBufferIn_short( 398);
	dataBufferOut_short( 381) <= dataBufferIn_short( 399);
	dataBufferOut_short( 464) <= dataBufferIn_short( 400);
	dataBufferOut_short( 547) <= dataBufferIn_short( 401);
	dataBufferOut_short( 630) <= dataBufferIn_short( 402);
	dataBufferOut_short( 713) <= dataBufferIn_short( 403);
	dataBufferOut_short( 796) <= dataBufferIn_short( 404);
	dataBufferOut_short( 879) <= dataBufferIn_short( 405);
	dataBufferOut_short( 962) <= dataBufferIn_short( 406);
	dataBufferOut_short(1045) <= dataBufferIn_short( 407);
	dataBufferOut_short(  72) <= dataBufferIn_short( 408);
	dataBufferOut_short( 155) <= dataBufferIn_short( 409);
	dataBufferOut_short( 238) <= dataBufferIn_short( 410);
	dataBufferOut_short( 321) <= dataBufferIn_short( 411);
	dataBufferOut_short( 404) <= dataBufferIn_short( 412);
	dataBufferOut_short( 487) <= dataBufferIn_short( 413);
	dataBufferOut_short( 570) <= dataBufferIn_short( 414);
	dataBufferOut_short( 653) <= dataBufferIn_short( 415);
	dataBufferOut_short( 736) <= dataBufferIn_short( 416);
	dataBufferOut_short( 819) <= dataBufferIn_short( 417);
	dataBufferOut_short( 902) <= dataBufferIn_short( 418);
	dataBufferOut_short( 985) <= dataBufferIn_short( 419);
	dataBufferOut_short(  12) <= dataBufferIn_short( 420);
	dataBufferOut_short(  95) <= dataBufferIn_short( 421);
	dataBufferOut_short( 178) <= dataBufferIn_short( 422);
	dataBufferOut_short( 261) <= dataBufferIn_short( 423);
	dataBufferOut_short( 344) <= dataBufferIn_short( 424);
	dataBufferOut_short( 427) <= dataBufferIn_short( 425);
	dataBufferOut_short( 510) <= dataBufferIn_short( 426);
	dataBufferOut_short( 593) <= dataBufferIn_short( 427);
	dataBufferOut_short( 676) <= dataBufferIn_short( 428);
	dataBufferOut_short( 759) <= dataBufferIn_short( 429);
	dataBufferOut_short( 842) <= dataBufferIn_short( 430);
	dataBufferOut_short( 925) <= dataBufferIn_short( 431);
	dataBufferOut_short(1008) <= dataBufferIn_short( 432);
	dataBufferOut_short(  35) <= dataBufferIn_short( 433);
	dataBufferOut_short( 118) <= dataBufferIn_short( 434);
	dataBufferOut_short( 201) <= dataBufferIn_short( 435);
	dataBufferOut_short( 284) <= dataBufferIn_short( 436);
	dataBufferOut_short( 367) <= dataBufferIn_short( 437);
	dataBufferOut_short( 450) <= dataBufferIn_short( 438);
	dataBufferOut_short( 533) <= dataBufferIn_short( 439);
	dataBufferOut_short( 616) <= dataBufferIn_short( 440);
	dataBufferOut_short( 699) <= dataBufferIn_short( 441);
	dataBufferOut_short( 782) <= dataBufferIn_short( 442);
	dataBufferOut_short( 865) <= dataBufferIn_short( 443);
	dataBufferOut_short( 948) <= dataBufferIn_short( 444);
	dataBufferOut_short(1031) <= dataBufferIn_short( 445);
	dataBufferOut_short(  58) <= dataBufferIn_short( 446);
	dataBufferOut_short( 141) <= dataBufferIn_short( 447);
	dataBufferOut_short( 224) <= dataBufferIn_short( 448);
	dataBufferOut_short( 307) <= dataBufferIn_short( 449);
	dataBufferOut_short( 390) <= dataBufferIn_short( 450);
	dataBufferOut_short( 473) <= dataBufferIn_short( 451);
	dataBufferOut_short( 556) <= dataBufferIn_short( 452);
	dataBufferOut_short( 639) <= dataBufferIn_short( 453);
	dataBufferOut_short( 722) <= dataBufferIn_short( 454);
	dataBufferOut_short( 805) <= dataBufferIn_short( 455);
	dataBufferOut_short( 888) <= dataBufferIn_short( 456);
	dataBufferOut_short( 971) <= dataBufferIn_short( 457);
	dataBufferOut_short(1054) <= dataBufferIn_short( 458);
	dataBufferOut_short(  81) <= dataBufferIn_short( 459);
	dataBufferOut_short( 164) <= dataBufferIn_short( 460);
	dataBufferOut_short( 247) <= dataBufferIn_short( 461);
	dataBufferOut_short( 330) <= dataBufferIn_short( 462);
	dataBufferOut_short( 413) <= dataBufferIn_short( 463);
	dataBufferOut_short( 496) <= dataBufferIn_short( 464);
	dataBufferOut_short( 579) <= dataBufferIn_short( 465);
	dataBufferOut_short( 662) <= dataBufferIn_short( 466);
	dataBufferOut_short( 745) <= dataBufferIn_short( 467);
	dataBufferOut_short( 828) <= dataBufferIn_short( 468);
	dataBufferOut_short( 911) <= dataBufferIn_short( 469);
	dataBufferOut_short( 994) <= dataBufferIn_short( 470);
	dataBufferOut_short(  21) <= dataBufferIn_short( 471);
	dataBufferOut_short( 104) <= dataBufferIn_short( 472);
	dataBufferOut_short( 187) <= dataBufferIn_short( 473);
	dataBufferOut_short( 270) <= dataBufferIn_short( 474);
	dataBufferOut_short( 353) <= dataBufferIn_short( 475);
	dataBufferOut_short( 436) <= dataBufferIn_short( 476);
	dataBufferOut_short( 519) <= dataBufferIn_short( 477);
	dataBufferOut_short( 602) <= dataBufferIn_short( 478);
	dataBufferOut_short( 685) <= dataBufferIn_short( 479);
	dataBufferOut_short( 768) <= dataBufferIn_short( 480);
	dataBufferOut_short( 851) <= dataBufferIn_short( 481);
	dataBufferOut_short( 934) <= dataBufferIn_short( 482);
	dataBufferOut_short(1017) <= dataBufferIn_short( 483);
	dataBufferOut_short(  44) <= dataBufferIn_short( 484);
	dataBufferOut_short( 127) <= dataBufferIn_short( 485);
	dataBufferOut_short( 210) <= dataBufferIn_short( 486);
	dataBufferOut_short( 293) <= dataBufferIn_short( 487);
	dataBufferOut_short( 376) <= dataBufferIn_short( 488);
	dataBufferOut_short( 459) <= dataBufferIn_short( 489);
	dataBufferOut_short( 542) <= dataBufferIn_short( 490);
	dataBufferOut_short( 625) <= dataBufferIn_short( 491);
	dataBufferOut_short( 708) <= dataBufferIn_short( 492);
	dataBufferOut_short( 791) <= dataBufferIn_short( 493);
	dataBufferOut_short( 874) <= dataBufferIn_short( 494);
	dataBufferOut_short( 957) <= dataBufferIn_short( 495);
	dataBufferOut_short(1040) <= dataBufferIn_short( 496);
	dataBufferOut_short(  67) <= dataBufferIn_short( 497);
	dataBufferOut_short( 150) <= dataBufferIn_short( 498);
	dataBufferOut_short( 233) <= dataBufferIn_short( 499);
	dataBufferOut_short( 316) <= dataBufferIn_short( 500);
	dataBufferOut_short( 399) <= dataBufferIn_short( 501);
	dataBufferOut_short( 482) <= dataBufferIn_short( 502);
	dataBufferOut_short( 565) <= dataBufferIn_short( 503);
	dataBufferOut_short( 648) <= dataBufferIn_short( 504);
	dataBufferOut_short( 731) <= dataBufferIn_short( 505);
	dataBufferOut_short( 814) <= dataBufferIn_short( 506);
	dataBufferOut_short( 897) <= dataBufferIn_short( 507);
	dataBufferOut_short( 980) <= dataBufferIn_short( 508);
	dataBufferOut_short(   7) <= dataBufferIn_short( 509);
	dataBufferOut_short(  90) <= dataBufferIn_short( 510);
	dataBufferOut_short( 173) <= dataBufferIn_short( 511);
	dataBufferOut_short( 256) <= dataBufferIn_short( 512);
	dataBufferOut_short( 339) <= dataBufferIn_short( 513);
	dataBufferOut_short( 422) <= dataBufferIn_short( 514);
	dataBufferOut_short( 505) <= dataBufferIn_short( 515);
	dataBufferOut_short( 588) <= dataBufferIn_short( 516);
	dataBufferOut_short( 671) <= dataBufferIn_short( 517);
	dataBufferOut_short( 754) <= dataBufferIn_short( 518);
	dataBufferOut_short( 837) <= dataBufferIn_short( 519);
	dataBufferOut_short( 920) <= dataBufferIn_short( 520);
	dataBufferOut_short(1003) <= dataBufferIn_short( 521);
	dataBufferOut_short(  30) <= dataBufferIn_short( 522);
	dataBufferOut_short( 113) <= dataBufferIn_short( 523);
	dataBufferOut_short( 196) <= dataBufferIn_short( 524);
	dataBufferOut_short( 279) <= dataBufferIn_short( 525);
	dataBufferOut_short( 362) <= dataBufferIn_short( 526);
	dataBufferOut_short( 445) <= dataBufferIn_short( 527);
	dataBufferOut_short( 528) <= dataBufferIn_short( 528);
	dataBufferOut_short( 611) <= dataBufferIn_short( 529);
	dataBufferOut_short( 694) <= dataBufferIn_short( 530);
	dataBufferOut_short( 777) <= dataBufferIn_short( 531);
	dataBufferOut_short( 860) <= dataBufferIn_short( 532);
	dataBufferOut_short( 943) <= dataBufferIn_short( 533);
	dataBufferOut_short(1026) <= dataBufferIn_short( 534);
	dataBufferOut_short(  53) <= dataBufferIn_short( 535);
	dataBufferOut_short( 136) <= dataBufferIn_short( 536);
	dataBufferOut_short( 219) <= dataBufferIn_short( 537);
	dataBufferOut_short( 302) <= dataBufferIn_short( 538);
	dataBufferOut_short( 385) <= dataBufferIn_short( 539);
	dataBufferOut_short( 468) <= dataBufferIn_short( 540);
	dataBufferOut_short( 551) <= dataBufferIn_short( 541);
	dataBufferOut_short( 634) <= dataBufferIn_short( 542);
	dataBufferOut_short( 717) <= dataBufferIn_short( 543);
	dataBufferOut_short( 800) <= dataBufferIn_short( 544);
	dataBufferOut_short( 883) <= dataBufferIn_short( 545);
	dataBufferOut_short( 966) <= dataBufferIn_short( 546);
	dataBufferOut_short(1049) <= dataBufferIn_short( 547);
	dataBufferOut_short(  76) <= dataBufferIn_short( 548);
	dataBufferOut_short( 159) <= dataBufferIn_short( 549);
	dataBufferOut_short( 242) <= dataBufferIn_short( 550);
	dataBufferOut_short( 325) <= dataBufferIn_short( 551);
	dataBufferOut_short( 408) <= dataBufferIn_short( 552);
	dataBufferOut_short( 491) <= dataBufferIn_short( 553);
	dataBufferOut_short( 574) <= dataBufferIn_short( 554);
	dataBufferOut_short( 657) <= dataBufferIn_short( 555);
	dataBufferOut_short( 740) <= dataBufferIn_short( 556);
	dataBufferOut_short( 823) <= dataBufferIn_short( 557);
	dataBufferOut_short( 906) <= dataBufferIn_short( 558);
	dataBufferOut_short( 989) <= dataBufferIn_short( 559);
	dataBufferOut_short(  16) <= dataBufferIn_short( 560);
	dataBufferOut_short(  99) <= dataBufferIn_short( 561);
	dataBufferOut_short( 182) <= dataBufferIn_short( 562);
	dataBufferOut_short( 265) <= dataBufferIn_short( 563);
	dataBufferOut_short( 348) <= dataBufferIn_short( 564);
	dataBufferOut_short( 431) <= dataBufferIn_short( 565);
	dataBufferOut_short( 514) <= dataBufferIn_short( 566);
	dataBufferOut_short( 597) <= dataBufferIn_short( 567);
	dataBufferOut_short( 680) <= dataBufferIn_short( 568);
	dataBufferOut_short( 763) <= dataBufferIn_short( 569);
	dataBufferOut_short( 846) <= dataBufferIn_short( 570);
	dataBufferOut_short( 929) <= dataBufferIn_short( 571);
	dataBufferOut_short(1012) <= dataBufferIn_short( 572);
	dataBufferOut_short(  39) <= dataBufferIn_short( 573);
	dataBufferOut_short( 122) <= dataBufferIn_short( 574);
	dataBufferOut_short( 205) <= dataBufferIn_short( 575);
	dataBufferOut_short( 288) <= dataBufferIn_short( 576);
	dataBufferOut_short( 371) <= dataBufferIn_short( 577);
	dataBufferOut_short( 454) <= dataBufferIn_short( 578);
	dataBufferOut_short( 537) <= dataBufferIn_short( 579);
	dataBufferOut_short( 620) <= dataBufferIn_short( 580);
	dataBufferOut_short( 703) <= dataBufferIn_short( 581);
	dataBufferOut_short( 786) <= dataBufferIn_short( 582);
	dataBufferOut_short( 869) <= dataBufferIn_short( 583);
	dataBufferOut_short( 952) <= dataBufferIn_short( 584);
	dataBufferOut_short(1035) <= dataBufferIn_short( 585);
	dataBufferOut_short(  62) <= dataBufferIn_short( 586);
	dataBufferOut_short( 145) <= dataBufferIn_short( 587);
	dataBufferOut_short( 228) <= dataBufferIn_short( 588);
	dataBufferOut_short( 311) <= dataBufferIn_short( 589);
	dataBufferOut_short( 394) <= dataBufferIn_short( 590);
	dataBufferOut_short( 477) <= dataBufferIn_short( 591);
	dataBufferOut_short( 560) <= dataBufferIn_short( 592);
	dataBufferOut_short( 643) <= dataBufferIn_short( 593);
	dataBufferOut_short( 726) <= dataBufferIn_short( 594);
	dataBufferOut_short( 809) <= dataBufferIn_short( 595);
	dataBufferOut_short( 892) <= dataBufferIn_short( 596);
	dataBufferOut_short( 975) <= dataBufferIn_short( 597);
	dataBufferOut_short(   2) <= dataBufferIn_short( 598);
	dataBufferOut_short(  85) <= dataBufferIn_short( 599);
	dataBufferOut_short( 168) <= dataBufferIn_short( 600);
	dataBufferOut_short( 251) <= dataBufferIn_short( 601);
	dataBufferOut_short( 334) <= dataBufferIn_short( 602);
	dataBufferOut_short( 417) <= dataBufferIn_short( 603);
	dataBufferOut_short( 500) <= dataBufferIn_short( 604);
	dataBufferOut_short( 583) <= dataBufferIn_short( 605);
	dataBufferOut_short( 666) <= dataBufferIn_short( 606);
	dataBufferOut_short( 749) <= dataBufferIn_short( 607);
	dataBufferOut_short( 832) <= dataBufferIn_short( 608);
	dataBufferOut_short( 915) <= dataBufferIn_short( 609);
	dataBufferOut_short( 998) <= dataBufferIn_short( 610);
	dataBufferOut_short(  25) <= dataBufferIn_short( 611);
	dataBufferOut_short( 108) <= dataBufferIn_short( 612);
	dataBufferOut_short( 191) <= dataBufferIn_short( 613);
	dataBufferOut_short( 274) <= dataBufferIn_short( 614);
	dataBufferOut_short( 357) <= dataBufferIn_short( 615);
	dataBufferOut_short( 440) <= dataBufferIn_short( 616);
	dataBufferOut_short( 523) <= dataBufferIn_short( 617);
	dataBufferOut_short( 606) <= dataBufferIn_short( 618);
	dataBufferOut_short( 689) <= dataBufferIn_short( 619);
	dataBufferOut_short( 772) <= dataBufferIn_short( 620);
	dataBufferOut_short( 855) <= dataBufferIn_short( 621);
	dataBufferOut_short( 938) <= dataBufferIn_short( 622);
	dataBufferOut_short(1021) <= dataBufferIn_short( 623);
	dataBufferOut_short(  48) <= dataBufferIn_short( 624);
	dataBufferOut_short( 131) <= dataBufferIn_short( 625);
	dataBufferOut_short( 214) <= dataBufferIn_short( 626);
	dataBufferOut_short( 297) <= dataBufferIn_short( 627);
	dataBufferOut_short( 380) <= dataBufferIn_short( 628);
	dataBufferOut_short( 463) <= dataBufferIn_short( 629);
	dataBufferOut_short( 546) <= dataBufferIn_short( 630);
	dataBufferOut_short( 629) <= dataBufferIn_short( 631);
	dataBufferOut_short( 712) <= dataBufferIn_short( 632);
	dataBufferOut_short( 795) <= dataBufferIn_short( 633);
	dataBufferOut_short( 878) <= dataBufferIn_short( 634);
	dataBufferOut_short( 961) <= dataBufferIn_short( 635);
	dataBufferOut_short(1044) <= dataBufferIn_short( 636);
	dataBufferOut_short(  71) <= dataBufferIn_short( 637);
	dataBufferOut_short( 154) <= dataBufferIn_short( 638);
	dataBufferOut_short( 237) <= dataBufferIn_short( 639);
	dataBufferOut_short( 320) <= dataBufferIn_short( 640);
	dataBufferOut_short( 403) <= dataBufferIn_short( 641);
	dataBufferOut_short( 486) <= dataBufferIn_short( 642);
	dataBufferOut_short( 569) <= dataBufferIn_short( 643);
	dataBufferOut_short( 652) <= dataBufferIn_short( 644);
	dataBufferOut_short( 735) <= dataBufferIn_short( 645);
	dataBufferOut_short( 818) <= dataBufferIn_short( 646);
	dataBufferOut_short( 901) <= dataBufferIn_short( 647);
	dataBufferOut_short( 984) <= dataBufferIn_short( 648);
	dataBufferOut_short(  11) <= dataBufferIn_short( 649);
	dataBufferOut_short(  94) <= dataBufferIn_short( 650);
	dataBufferOut_short( 177) <= dataBufferIn_short( 651);
	dataBufferOut_short( 260) <= dataBufferIn_short( 652);
	dataBufferOut_short( 343) <= dataBufferIn_short( 653);
	dataBufferOut_short( 426) <= dataBufferIn_short( 654);
	dataBufferOut_short( 509) <= dataBufferIn_short( 655);
	dataBufferOut_short( 592) <= dataBufferIn_short( 656);
	dataBufferOut_short( 675) <= dataBufferIn_short( 657);
	dataBufferOut_short( 758) <= dataBufferIn_short( 658);
	dataBufferOut_short( 841) <= dataBufferIn_short( 659);
	dataBufferOut_short( 924) <= dataBufferIn_short( 660);
	dataBufferOut_short(1007) <= dataBufferIn_short( 661);
	dataBufferOut_short(  34) <= dataBufferIn_short( 662);
	dataBufferOut_short( 117) <= dataBufferIn_short( 663);
	dataBufferOut_short( 200) <= dataBufferIn_short( 664);
	dataBufferOut_short( 283) <= dataBufferIn_short( 665);
	dataBufferOut_short( 366) <= dataBufferIn_short( 666);
	dataBufferOut_short( 449) <= dataBufferIn_short( 667);
	dataBufferOut_short( 532) <= dataBufferIn_short( 668);
	dataBufferOut_short( 615) <= dataBufferIn_short( 669);
	dataBufferOut_short( 698) <= dataBufferIn_short( 670);
	dataBufferOut_short( 781) <= dataBufferIn_short( 671);
	dataBufferOut_short( 864) <= dataBufferIn_short( 672);
	dataBufferOut_short( 947) <= dataBufferIn_short( 673);
	dataBufferOut_short(1030) <= dataBufferIn_short( 674);
	dataBufferOut_short(  57) <= dataBufferIn_short( 675);
	dataBufferOut_short( 140) <= dataBufferIn_short( 676);
	dataBufferOut_short( 223) <= dataBufferIn_short( 677);
	dataBufferOut_short( 306) <= dataBufferIn_short( 678);
	dataBufferOut_short( 389) <= dataBufferIn_short( 679);
	dataBufferOut_short( 472) <= dataBufferIn_short( 680);
	dataBufferOut_short( 555) <= dataBufferIn_short( 681);
	dataBufferOut_short( 638) <= dataBufferIn_short( 682);
	dataBufferOut_short( 721) <= dataBufferIn_short( 683);
	dataBufferOut_short( 804) <= dataBufferIn_short( 684);
	dataBufferOut_short( 887) <= dataBufferIn_short( 685);
	dataBufferOut_short( 970) <= dataBufferIn_short( 686);
	dataBufferOut_short(1053) <= dataBufferIn_short( 687);
	dataBufferOut_short(  80) <= dataBufferIn_short( 688);
	dataBufferOut_short( 163) <= dataBufferIn_short( 689);
	dataBufferOut_short( 246) <= dataBufferIn_short( 690);
	dataBufferOut_short( 329) <= dataBufferIn_short( 691);
	dataBufferOut_short( 412) <= dataBufferIn_short( 692);
	dataBufferOut_short( 495) <= dataBufferIn_short( 693);
	dataBufferOut_short( 578) <= dataBufferIn_short( 694);
	dataBufferOut_short( 661) <= dataBufferIn_short( 695);
	dataBufferOut_short( 744) <= dataBufferIn_short( 696);
	dataBufferOut_short( 827) <= dataBufferIn_short( 697);
	dataBufferOut_short( 910) <= dataBufferIn_short( 698);
	dataBufferOut_short( 993) <= dataBufferIn_short( 699);
	dataBufferOut_short(  20) <= dataBufferIn_short( 700);
	dataBufferOut_short( 103) <= dataBufferIn_short( 701);
	dataBufferOut_short( 186) <= dataBufferIn_short( 702);
	dataBufferOut_short( 269) <= dataBufferIn_short( 703);
	dataBufferOut_short( 352) <= dataBufferIn_short( 704);
	dataBufferOut_short( 435) <= dataBufferIn_short( 705);
	dataBufferOut_short( 518) <= dataBufferIn_short( 706);
	dataBufferOut_short( 601) <= dataBufferIn_short( 707);
	dataBufferOut_short( 684) <= dataBufferIn_short( 708);
	dataBufferOut_short( 767) <= dataBufferIn_short( 709);
	dataBufferOut_short( 850) <= dataBufferIn_short( 710);
	dataBufferOut_short( 933) <= dataBufferIn_short( 711);
	dataBufferOut_short(1016) <= dataBufferIn_short( 712);
	dataBufferOut_short(  43) <= dataBufferIn_short( 713);
	dataBufferOut_short( 126) <= dataBufferIn_short( 714);
	dataBufferOut_short( 209) <= dataBufferIn_short( 715);
	dataBufferOut_short( 292) <= dataBufferIn_short( 716);
	dataBufferOut_short( 375) <= dataBufferIn_short( 717);
	dataBufferOut_short( 458) <= dataBufferIn_short( 718);
	dataBufferOut_short( 541) <= dataBufferIn_short( 719);
	dataBufferOut_short( 624) <= dataBufferIn_short( 720);
	dataBufferOut_short( 707) <= dataBufferIn_short( 721);
	dataBufferOut_short( 790) <= dataBufferIn_short( 722);
	dataBufferOut_short( 873) <= dataBufferIn_short( 723);
	dataBufferOut_short( 956) <= dataBufferIn_short( 724);
	dataBufferOut_short(1039) <= dataBufferIn_short( 725);
	dataBufferOut_short(  66) <= dataBufferIn_short( 726);
	dataBufferOut_short( 149) <= dataBufferIn_short( 727);
	dataBufferOut_short( 232) <= dataBufferIn_short( 728);
	dataBufferOut_short( 315) <= dataBufferIn_short( 729);
	dataBufferOut_short( 398) <= dataBufferIn_short( 730);
	dataBufferOut_short( 481) <= dataBufferIn_short( 731);
	dataBufferOut_short( 564) <= dataBufferIn_short( 732);
	dataBufferOut_short( 647) <= dataBufferIn_short( 733);
	dataBufferOut_short( 730) <= dataBufferIn_short( 734);
	dataBufferOut_short( 813) <= dataBufferIn_short( 735);
	dataBufferOut_short( 896) <= dataBufferIn_short( 736);
	dataBufferOut_short( 979) <= dataBufferIn_short( 737);
	dataBufferOut_short(   6) <= dataBufferIn_short( 738);
	dataBufferOut_short(  89) <= dataBufferIn_short( 739);
	dataBufferOut_short( 172) <= dataBufferIn_short( 740);
	dataBufferOut_short( 255) <= dataBufferIn_short( 741);
	dataBufferOut_short( 338) <= dataBufferIn_short( 742);
	dataBufferOut_short( 421) <= dataBufferIn_short( 743);
	dataBufferOut_short( 504) <= dataBufferIn_short( 744);
	dataBufferOut_short( 587) <= dataBufferIn_short( 745);
	dataBufferOut_short( 670) <= dataBufferIn_short( 746);
	dataBufferOut_short( 753) <= dataBufferIn_short( 747);
	dataBufferOut_short( 836) <= dataBufferIn_short( 748);
	dataBufferOut_short( 919) <= dataBufferIn_short( 749);
	dataBufferOut_short(1002) <= dataBufferIn_short( 750);
	dataBufferOut_short(  29) <= dataBufferIn_short( 751);
	dataBufferOut_short( 112) <= dataBufferIn_short( 752);
	dataBufferOut_short( 195) <= dataBufferIn_short( 753);
	dataBufferOut_short( 278) <= dataBufferIn_short( 754);
	dataBufferOut_short( 361) <= dataBufferIn_short( 755);
	dataBufferOut_short( 444) <= dataBufferIn_short( 756);
	dataBufferOut_short( 527) <= dataBufferIn_short( 757);
	dataBufferOut_short( 610) <= dataBufferIn_short( 758);
	dataBufferOut_short( 693) <= dataBufferIn_short( 759);
	dataBufferOut_short( 776) <= dataBufferIn_short( 760);
	dataBufferOut_short( 859) <= dataBufferIn_short( 761);
	dataBufferOut_short( 942) <= dataBufferIn_short( 762);
	dataBufferOut_short(1025) <= dataBufferIn_short( 763);
	dataBufferOut_short(  52) <= dataBufferIn_short( 764);
	dataBufferOut_short( 135) <= dataBufferIn_short( 765);
	dataBufferOut_short( 218) <= dataBufferIn_short( 766);
	dataBufferOut_short( 301) <= dataBufferIn_short( 767);
	dataBufferOut_short( 384) <= dataBufferIn_short( 768);
	dataBufferOut_short( 467) <= dataBufferIn_short( 769);
	dataBufferOut_short( 550) <= dataBufferIn_short( 770);
	dataBufferOut_short( 633) <= dataBufferIn_short( 771);
	dataBufferOut_short( 716) <= dataBufferIn_short( 772);
	dataBufferOut_short( 799) <= dataBufferIn_short( 773);
	dataBufferOut_short( 882) <= dataBufferIn_short( 774);
	dataBufferOut_short( 965) <= dataBufferIn_short( 775);
	dataBufferOut_short(1048) <= dataBufferIn_short( 776);
	dataBufferOut_short(  75) <= dataBufferIn_short( 777);
	dataBufferOut_short( 158) <= dataBufferIn_short( 778);
	dataBufferOut_short( 241) <= dataBufferIn_short( 779);
	dataBufferOut_short( 324) <= dataBufferIn_short( 780);
	dataBufferOut_short( 407) <= dataBufferIn_short( 781);
	dataBufferOut_short( 490) <= dataBufferIn_short( 782);
	dataBufferOut_short( 573) <= dataBufferIn_short( 783);
	dataBufferOut_short( 656) <= dataBufferIn_short( 784);
	dataBufferOut_short( 739) <= dataBufferIn_short( 785);
	dataBufferOut_short( 822) <= dataBufferIn_short( 786);
	dataBufferOut_short( 905) <= dataBufferIn_short( 787);
	dataBufferOut_short( 988) <= dataBufferIn_short( 788);
	dataBufferOut_short(  15) <= dataBufferIn_short( 789);
	dataBufferOut_short(  98) <= dataBufferIn_short( 790);
	dataBufferOut_short( 181) <= dataBufferIn_short( 791);
	dataBufferOut_short( 264) <= dataBufferIn_short( 792);
	dataBufferOut_short( 347) <= dataBufferIn_short( 793);
	dataBufferOut_short( 430) <= dataBufferIn_short( 794);
	dataBufferOut_short( 513) <= dataBufferIn_short( 795);
	dataBufferOut_short( 596) <= dataBufferIn_short( 796);
	dataBufferOut_short( 679) <= dataBufferIn_short( 797);
	dataBufferOut_short( 762) <= dataBufferIn_short( 798);
	dataBufferOut_short( 845) <= dataBufferIn_short( 799);
	dataBufferOut_short( 928) <= dataBufferIn_short( 800);
	dataBufferOut_short(1011) <= dataBufferIn_short( 801);
	dataBufferOut_short(  38) <= dataBufferIn_short( 802);
	dataBufferOut_short( 121) <= dataBufferIn_short( 803);
	dataBufferOut_short( 204) <= dataBufferIn_short( 804);
	dataBufferOut_short( 287) <= dataBufferIn_short( 805);
	dataBufferOut_short( 370) <= dataBufferIn_short( 806);
	dataBufferOut_short( 453) <= dataBufferIn_short( 807);
	dataBufferOut_short( 536) <= dataBufferIn_short( 808);
	dataBufferOut_short( 619) <= dataBufferIn_short( 809);
	dataBufferOut_short( 702) <= dataBufferIn_short( 810);
	dataBufferOut_short( 785) <= dataBufferIn_short( 811);
	dataBufferOut_short( 868) <= dataBufferIn_short( 812);
	dataBufferOut_short( 951) <= dataBufferIn_short( 813);
	dataBufferOut_short(1034) <= dataBufferIn_short( 814);
	dataBufferOut_short(  61) <= dataBufferIn_short( 815);
	dataBufferOut_short( 144) <= dataBufferIn_short( 816);
	dataBufferOut_short( 227) <= dataBufferIn_short( 817);
	dataBufferOut_short( 310) <= dataBufferIn_short( 818);
	dataBufferOut_short( 393) <= dataBufferIn_short( 819);
	dataBufferOut_short( 476) <= dataBufferIn_short( 820);
	dataBufferOut_short( 559) <= dataBufferIn_short( 821);
	dataBufferOut_short( 642) <= dataBufferIn_short( 822);
	dataBufferOut_short( 725) <= dataBufferIn_short( 823);
	dataBufferOut_short( 808) <= dataBufferIn_short( 824);
	dataBufferOut_short( 891) <= dataBufferIn_short( 825);
	dataBufferOut_short( 974) <= dataBufferIn_short( 826);
	dataBufferOut_short(   1) <= dataBufferIn_short( 827);
	dataBufferOut_short(  84) <= dataBufferIn_short( 828);
	dataBufferOut_short( 167) <= dataBufferIn_short( 829);
	dataBufferOut_short( 250) <= dataBufferIn_short( 830);
	dataBufferOut_short( 333) <= dataBufferIn_short( 831);
	dataBufferOut_short( 416) <= dataBufferIn_short( 832);
	dataBufferOut_short( 499) <= dataBufferIn_short( 833);
	dataBufferOut_short( 582) <= dataBufferIn_short( 834);
	dataBufferOut_short( 665) <= dataBufferIn_short( 835);
	dataBufferOut_short( 748) <= dataBufferIn_short( 836);
	dataBufferOut_short( 831) <= dataBufferIn_short( 837);
	dataBufferOut_short( 914) <= dataBufferIn_short( 838);
	dataBufferOut_short( 997) <= dataBufferIn_short( 839);
	dataBufferOut_short(  24) <= dataBufferIn_short( 840);
	dataBufferOut_short( 107) <= dataBufferIn_short( 841);
	dataBufferOut_short( 190) <= dataBufferIn_short( 842);
	dataBufferOut_short( 273) <= dataBufferIn_short( 843);
	dataBufferOut_short( 356) <= dataBufferIn_short( 844);
	dataBufferOut_short( 439) <= dataBufferIn_short( 845);
	dataBufferOut_short( 522) <= dataBufferIn_short( 846);
	dataBufferOut_short( 605) <= dataBufferIn_short( 847);
	dataBufferOut_short( 688) <= dataBufferIn_short( 848);
	dataBufferOut_short( 771) <= dataBufferIn_short( 849);
	dataBufferOut_short( 854) <= dataBufferIn_short( 850);
	dataBufferOut_short( 937) <= dataBufferIn_short( 851);
	dataBufferOut_short(1020) <= dataBufferIn_short( 852);
	dataBufferOut_short(  47) <= dataBufferIn_short( 853);
	dataBufferOut_short( 130) <= dataBufferIn_short( 854);
	dataBufferOut_short( 213) <= dataBufferIn_short( 855);
	dataBufferOut_short( 296) <= dataBufferIn_short( 856);
	dataBufferOut_short( 379) <= dataBufferIn_short( 857);
	dataBufferOut_short( 462) <= dataBufferIn_short( 858);
	dataBufferOut_short( 545) <= dataBufferIn_short( 859);
	dataBufferOut_short( 628) <= dataBufferIn_short( 860);
	dataBufferOut_short( 711) <= dataBufferIn_short( 861);
	dataBufferOut_short( 794) <= dataBufferIn_short( 862);
	dataBufferOut_short( 877) <= dataBufferIn_short( 863);
	dataBufferOut_short( 960) <= dataBufferIn_short( 864);
	dataBufferOut_short(1043) <= dataBufferIn_short( 865);
	dataBufferOut_short(  70) <= dataBufferIn_short( 866);
	dataBufferOut_short( 153) <= dataBufferIn_short( 867);
	dataBufferOut_short( 236) <= dataBufferIn_short( 868);
	dataBufferOut_short( 319) <= dataBufferIn_short( 869);
	dataBufferOut_short( 402) <= dataBufferIn_short( 870);
	dataBufferOut_short( 485) <= dataBufferIn_short( 871);
	dataBufferOut_short( 568) <= dataBufferIn_short( 872);
	dataBufferOut_short( 651) <= dataBufferIn_short( 873);
	dataBufferOut_short( 734) <= dataBufferIn_short( 874);
	dataBufferOut_short( 817) <= dataBufferIn_short( 875);
	dataBufferOut_short( 900) <= dataBufferIn_short( 876);
	dataBufferOut_short( 983) <= dataBufferIn_short( 877);
	dataBufferOut_short(  10) <= dataBufferIn_short( 878);
	dataBufferOut_short(  93) <= dataBufferIn_short( 879);
	dataBufferOut_short( 176) <= dataBufferIn_short( 880);
	dataBufferOut_short( 259) <= dataBufferIn_short( 881);
	dataBufferOut_short( 342) <= dataBufferIn_short( 882);
	dataBufferOut_short( 425) <= dataBufferIn_short( 883);
	dataBufferOut_short( 508) <= dataBufferIn_short( 884);
	dataBufferOut_short( 591) <= dataBufferIn_short( 885);
	dataBufferOut_short( 674) <= dataBufferIn_short( 886);
	dataBufferOut_short( 757) <= dataBufferIn_short( 887);
	dataBufferOut_short( 840) <= dataBufferIn_short( 888);
	dataBufferOut_short( 923) <= dataBufferIn_short( 889);
	dataBufferOut_short(1006) <= dataBufferIn_short( 890);
	dataBufferOut_short(  33) <= dataBufferIn_short( 891);
	dataBufferOut_short( 116) <= dataBufferIn_short( 892);
	dataBufferOut_short( 199) <= dataBufferIn_short( 893);
	dataBufferOut_short( 282) <= dataBufferIn_short( 894);
	dataBufferOut_short( 365) <= dataBufferIn_short( 895);
	dataBufferOut_short( 448) <= dataBufferIn_short( 896);
	dataBufferOut_short( 531) <= dataBufferIn_short( 897);
	dataBufferOut_short( 614) <= dataBufferIn_short( 898);
	dataBufferOut_short( 697) <= dataBufferIn_short( 899);
	dataBufferOut_short( 780) <= dataBufferIn_short( 900);
	dataBufferOut_short( 863) <= dataBufferIn_short( 901);
	dataBufferOut_short( 946) <= dataBufferIn_short( 902);
	dataBufferOut_short(1029) <= dataBufferIn_short( 903);
	dataBufferOut_short(  56) <= dataBufferIn_short( 904);
	dataBufferOut_short( 139) <= dataBufferIn_short( 905);
	dataBufferOut_short( 222) <= dataBufferIn_short( 906);
	dataBufferOut_short( 305) <= dataBufferIn_short( 907);
	dataBufferOut_short( 388) <= dataBufferIn_short( 908);
	dataBufferOut_short( 471) <= dataBufferIn_short( 909);
	dataBufferOut_short( 554) <= dataBufferIn_short( 910);
	dataBufferOut_short( 637) <= dataBufferIn_short( 911);
	dataBufferOut_short( 720) <= dataBufferIn_short( 912);
	dataBufferOut_short( 803) <= dataBufferIn_short( 913);
	dataBufferOut_short( 886) <= dataBufferIn_short( 914);
	dataBufferOut_short( 969) <= dataBufferIn_short( 915);
	dataBufferOut_short(1052) <= dataBufferIn_short( 916);
	dataBufferOut_short(  79) <= dataBufferIn_short( 917);
	dataBufferOut_short( 162) <= dataBufferIn_short( 918);
	dataBufferOut_short( 245) <= dataBufferIn_short( 919);
	dataBufferOut_short( 328) <= dataBufferIn_short( 920);
	dataBufferOut_short( 411) <= dataBufferIn_short( 921);
	dataBufferOut_short( 494) <= dataBufferIn_short( 922);
	dataBufferOut_short( 577) <= dataBufferIn_short( 923);
	dataBufferOut_short( 660) <= dataBufferIn_short( 924);
	dataBufferOut_short( 743) <= dataBufferIn_short( 925);
	dataBufferOut_short( 826) <= dataBufferIn_short( 926);
	dataBufferOut_short( 909) <= dataBufferIn_short( 927);
	dataBufferOut_short( 992) <= dataBufferIn_short( 928);
	dataBufferOut_short(  19) <= dataBufferIn_short( 929);
	dataBufferOut_short( 102) <= dataBufferIn_short( 930);
	dataBufferOut_short( 185) <= dataBufferIn_short( 931);
	dataBufferOut_short( 268) <= dataBufferIn_short( 932);
	dataBufferOut_short( 351) <= dataBufferIn_short( 933);
	dataBufferOut_short( 434) <= dataBufferIn_short( 934);
	dataBufferOut_short( 517) <= dataBufferIn_short( 935);
	dataBufferOut_short( 600) <= dataBufferIn_short( 936);
	dataBufferOut_short( 683) <= dataBufferIn_short( 937);
	dataBufferOut_short( 766) <= dataBufferIn_short( 938);
	dataBufferOut_short( 849) <= dataBufferIn_short( 939);
	dataBufferOut_short( 932) <= dataBufferIn_short( 940);
	dataBufferOut_short(1015) <= dataBufferIn_short( 941);
	dataBufferOut_short(  42) <= dataBufferIn_short( 942);
	dataBufferOut_short( 125) <= dataBufferIn_short( 943);
	dataBufferOut_short( 208) <= dataBufferIn_short( 944);
	dataBufferOut_short( 291) <= dataBufferIn_short( 945);
	dataBufferOut_short( 374) <= dataBufferIn_short( 946);
	dataBufferOut_short( 457) <= dataBufferIn_short( 947);
	dataBufferOut_short( 540) <= dataBufferIn_short( 948);
	dataBufferOut_short( 623) <= dataBufferIn_short( 949);
	dataBufferOut_short( 706) <= dataBufferIn_short( 950);
	dataBufferOut_short( 789) <= dataBufferIn_short( 951);
	dataBufferOut_short( 872) <= dataBufferIn_short( 952);
	dataBufferOut_short( 955) <= dataBufferIn_short( 953);
	dataBufferOut_short(1038) <= dataBufferIn_short( 954);
	dataBufferOut_short(  65) <= dataBufferIn_short( 955);
	dataBufferOut_short( 148) <= dataBufferIn_short( 956);
	dataBufferOut_short( 231) <= dataBufferIn_short( 957);
	dataBufferOut_short( 314) <= dataBufferIn_short( 958);
	dataBufferOut_short( 397) <= dataBufferIn_short( 959);
	dataBufferOut_short( 480) <= dataBufferIn_short( 960);
	dataBufferOut_short( 563) <= dataBufferIn_short( 961);
	dataBufferOut_short( 646) <= dataBufferIn_short( 962);
	dataBufferOut_short( 729) <= dataBufferIn_short( 963);
	dataBufferOut_short( 812) <= dataBufferIn_short( 964);
	dataBufferOut_short( 895) <= dataBufferIn_short( 965);
	dataBufferOut_short( 978) <= dataBufferIn_short( 966);
	dataBufferOut_short(   5) <= dataBufferIn_short( 967);
	dataBufferOut_short(  88) <= dataBufferIn_short( 968);
	dataBufferOut_short( 171) <= dataBufferIn_short( 969);
	dataBufferOut_short( 254) <= dataBufferIn_short( 970);
	dataBufferOut_short( 337) <= dataBufferIn_short( 971);
	dataBufferOut_short( 420) <= dataBufferIn_short( 972);
	dataBufferOut_short( 503) <= dataBufferIn_short( 973);
	dataBufferOut_short( 586) <= dataBufferIn_short( 974);
	dataBufferOut_short( 669) <= dataBufferIn_short( 975);
	dataBufferOut_short( 752) <= dataBufferIn_short( 976);
	dataBufferOut_short( 835) <= dataBufferIn_short( 977);
	dataBufferOut_short( 918) <= dataBufferIn_short( 978);
	dataBufferOut_short(1001) <= dataBufferIn_short( 979);
	dataBufferOut_short(  28) <= dataBufferIn_short( 980);
	dataBufferOut_short( 111) <= dataBufferIn_short( 981);
	dataBufferOut_short( 194) <= dataBufferIn_short( 982);
	dataBufferOut_short( 277) <= dataBufferIn_short( 983);
	dataBufferOut_short( 360) <= dataBufferIn_short( 984);
	dataBufferOut_short( 443) <= dataBufferIn_short( 985);
	dataBufferOut_short( 526) <= dataBufferIn_short( 986);
	dataBufferOut_short( 609) <= dataBufferIn_short( 987);
	dataBufferOut_short( 692) <= dataBufferIn_short( 988);
	dataBufferOut_short( 775) <= dataBufferIn_short( 989);
	dataBufferOut_short( 858) <= dataBufferIn_short( 990);
	dataBufferOut_short( 941) <= dataBufferIn_short( 991);
	dataBufferOut_short(1024) <= dataBufferIn_short( 992);
	dataBufferOut_short(  51) <= dataBufferIn_short( 993);
	dataBufferOut_short( 134) <= dataBufferIn_short( 994);
	dataBufferOut_short( 217) <= dataBufferIn_short( 995);
	dataBufferOut_short( 300) <= dataBufferIn_short( 996);
	dataBufferOut_short( 383) <= dataBufferIn_short( 997);
	dataBufferOut_short( 466) <= dataBufferIn_short( 998);
	dataBufferOut_short( 549) <= dataBufferIn_short( 999);
	dataBufferOut_short( 632) <= dataBufferIn_short(1000);
	dataBufferOut_short( 715) <= dataBufferIn_short(1001);
	dataBufferOut_short( 798) <= dataBufferIn_short(1002);
	dataBufferOut_short( 881) <= dataBufferIn_short(1003);
	dataBufferOut_short( 964) <= dataBufferIn_short(1004);
	dataBufferOut_short(1047) <= dataBufferIn_short(1005);
	dataBufferOut_short(  74) <= dataBufferIn_short(1006);
	dataBufferOut_short( 157) <= dataBufferIn_short(1007);
	dataBufferOut_short( 240) <= dataBufferIn_short(1008);
	dataBufferOut_short( 323) <= dataBufferIn_short(1009);
	dataBufferOut_short( 406) <= dataBufferIn_short(1010);
	dataBufferOut_short( 489) <= dataBufferIn_short(1011);
	dataBufferOut_short( 572) <= dataBufferIn_short(1012);
	dataBufferOut_short( 655) <= dataBufferIn_short(1013);
	dataBufferOut_short( 738) <= dataBufferIn_short(1014);
	dataBufferOut_short( 821) <= dataBufferIn_short(1015);
	dataBufferOut_short( 904) <= dataBufferIn_short(1016);
	dataBufferOut_short( 987) <= dataBufferIn_short(1017);
	dataBufferOut_short(  14) <= dataBufferIn_short(1018);
	dataBufferOut_short(  97) <= dataBufferIn_short(1019);
	dataBufferOut_short( 180) <= dataBufferIn_short(1020);
	dataBufferOut_short( 263) <= dataBufferIn_short(1021);
	dataBufferOut_short( 346) <= dataBufferIn_short(1022);
	dataBufferOut_short( 429) <= dataBufferIn_short(1023);
	dataBufferOut_short( 512) <= dataBufferIn_short(1024);
	dataBufferOut_short( 595) <= dataBufferIn_short(1025);
	dataBufferOut_short( 678) <= dataBufferIn_short(1026);
	dataBufferOut_short( 761) <= dataBufferIn_short(1027);
	dataBufferOut_short( 844) <= dataBufferIn_short(1028);
	dataBufferOut_short( 927) <= dataBufferIn_short(1029);
	dataBufferOut_short(1010) <= dataBufferIn_short(1030);
	dataBufferOut_short(  37) <= dataBufferIn_short(1031);
	dataBufferOut_short( 120) <= dataBufferIn_short(1032);
	dataBufferOut_short( 203) <= dataBufferIn_short(1033);
	dataBufferOut_short( 286) <= dataBufferIn_short(1034);
	dataBufferOut_short( 369) <= dataBufferIn_short(1035);
	dataBufferOut_short( 452) <= dataBufferIn_short(1036);
	dataBufferOut_short( 535) <= dataBufferIn_short(1037);
	dataBufferOut_short( 618) <= dataBufferIn_short(1038);
	dataBufferOut_short( 701) <= dataBufferIn_short(1039);
	dataBufferOut_short( 784) <= dataBufferIn_short(1040);
	dataBufferOut_short( 867) <= dataBufferIn_short(1041);
	dataBufferOut_short( 950) <= dataBufferIn_short(1042);
	dataBufferOut_short(1033) <= dataBufferIn_short(1043);
	dataBufferOut_short(  60) <= dataBufferIn_short(1044);
	dataBufferOut_short( 143) <= dataBufferIn_short(1045);
	dataBufferOut_short( 226) <= dataBufferIn_short(1046);
	dataBufferOut_short( 309) <= dataBufferIn_short(1047);
	dataBufferOut_short( 392) <= dataBufferIn_short(1048);
	dataBufferOut_short( 475) <= dataBufferIn_short(1049);
	dataBufferOut_short( 558) <= dataBufferIn_short(1050);
	dataBufferOut_short( 641) <= dataBufferIn_short(1051);
	dataBufferOut_short( 724) <= dataBufferIn_short(1052);
	dataBufferOut_short( 807) <= dataBufferIn_short(1053);
	dataBufferOut_short( 890) <= dataBufferIn_short(1054);
	dataBufferOut_short( 973) <= dataBufferIn_short(1055);
	dataBufferOut_long(   0) <= dataBufferIn_long(   0);
	dataBufferOut_long( 743) <= dataBufferIn_long(   1);
	dataBufferOut_long(1486) <= dataBufferIn_long(   2);
	dataBufferOut_long(2229) <= dataBufferIn_long(   3);
	dataBufferOut_long(2972) <= dataBufferIn_long(   4);
	dataBufferOut_long(3715) <= dataBufferIn_long(   5);
	dataBufferOut_long(4458) <= dataBufferIn_long(   6);
	dataBufferOut_long(5201) <= dataBufferIn_long(   7);
	dataBufferOut_long(5944) <= dataBufferIn_long(   8);
	dataBufferOut_long( 543) <= dataBufferIn_long(   9);
	dataBufferOut_long(1286) <= dataBufferIn_long(  10);
	dataBufferOut_long(2029) <= dataBufferIn_long(  11);
	dataBufferOut_long(2772) <= dataBufferIn_long(  12);
	dataBufferOut_long(3515) <= dataBufferIn_long(  13);
	dataBufferOut_long(4258) <= dataBufferIn_long(  14);
	dataBufferOut_long(5001) <= dataBufferIn_long(  15);
	dataBufferOut_long(5744) <= dataBufferIn_long(  16);
	dataBufferOut_long( 343) <= dataBufferIn_long(  17);
	dataBufferOut_long(1086) <= dataBufferIn_long(  18);
	dataBufferOut_long(1829) <= dataBufferIn_long(  19);
	dataBufferOut_long(2572) <= dataBufferIn_long(  20);
	dataBufferOut_long(3315) <= dataBufferIn_long(  21);
	dataBufferOut_long(4058) <= dataBufferIn_long(  22);
	dataBufferOut_long(4801) <= dataBufferIn_long(  23);
	dataBufferOut_long(5544) <= dataBufferIn_long(  24);
	dataBufferOut_long( 143) <= dataBufferIn_long(  25);
	dataBufferOut_long( 886) <= dataBufferIn_long(  26);
	dataBufferOut_long(1629) <= dataBufferIn_long(  27);
	dataBufferOut_long(2372) <= dataBufferIn_long(  28);
	dataBufferOut_long(3115) <= dataBufferIn_long(  29);
	dataBufferOut_long(3858) <= dataBufferIn_long(  30);
	dataBufferOut_long(4601) <= dataBufferIn_long(  31);
	dataBufferOut_long(5344) <= dataBufferIn_long(  32);
	dataBufferOut_long(6087) <= dataBufferIn_long(  33);
	dataBufferOut_long( 686) <= dataBufferIn_long(  34);
	dataBufferOut_long(1429) <= dataBufferIn_long(  35);
	dataBufferOut_long(2172) <= dataBufferIn_long(  36);
	dataBufferOut_long(2915) <= dataBufferIn_long(  37);
	dataBufferOut_long(3658) <= dataBufferIn_long(  38);
	dataBufferOut_long(4401) <= dataBufferIn_long(  39);
	dataBufferOut_long(5144) <= dataBufferIn_long(  40);
	dataBufferOut_long(5887) <= dataBufferIn_long(  41);
	dataBufferOut_long( 486) <= dataBufferIn_long(  42);
	dataBufferOut_long(1229) <= dataBufferIn_long(  43);
	dataBufferOut_long(1972) <= dataBufferIn_long(  44);
	dataBufferOut_long(2715) <= dataBufferIn_long(  45);
	dataBufferOut_long(3458) <= dataBufferIn_long(  46);
	dataBufferOut_long(4201) <= dataBufferIn_long(  47);
	dataBufferOut_long(4944) <= dataBufferIn_long(  48);
	dataBufferOut_long(5687) <= dataBufferIn_long(  49);
	dataBufferOut_long( 286) <= dataBufferIn_long(  50);
	dataBufferOut_long(1029) <= dataBufferIn_long(  51);
	dataBufferOut_long(1772) <= dataBufferIn_long(  52);
	dataBufferOut_long(2515) <= dataBufferIn_long(  53);
	dataBufferOut_long(3258) <= dataBufferIn_long(  54);
	dataBufferOut_long(4001) <= dataBufferIn_long(  55);
	dataBufferOut_long(4744) <= dataBufferIn_long(  56);
	dataBufferOut_long(5487) <= dataBufferIn_long(  57);
	dataBufferOut_long(  86) <= dataBufferIn_long(  58);
	dataBufferOut_long( 829) <= dataBufferIn_long(  59);
	dataBufferOut_long(1572) <= dataBufferIn_long(  60);
	dataBufferOut_long(2315) <= dataBufferIn_long(  61);
	dataBufferOut_long(3058) <= dataBufferIn_long(  62);
	dataBufferOut_long(3801) <= dataBufferIn_long(  63);
	dataBufferOut_long(4544) <= dataBufferIn_long(  64);
	dataBufferOut_long(5287) <= dataBufferIn_long(  65);
	dataBufferOut_long(6030) <= dataBufferIn_long(  66);
	dataBufferOut_long( 629) <= dataBufferIn_long(  67);
	dataBufferOut_long(1372) <= dataBufferIn_long(  68);
	dataBufferOut_long(2115) <= dataBufferIn_long(  69);
	dataBufferOut_long(2858) <= dataBufferIn_long(  70);
	dataBufferOut_long(3601) <= dataBufferIn_long(  71);
	dataBufferOut_long(4344) <= dataBufferIn_long(  72);
	dataBufferOut_long(5087) <= dataBufferIn_long(  73);
	dataBufferOut_long(5830) <= dataBufferIn_long(  74);
	dataBufferOut_long( 429) <= dataBufferIn_long(  75);
	dataBufferOut_long(1172) <= dataBufferIn_long(  76);
	dataBufferOut_long(1915) <= dataBufferIn_long(  77);
	dataBufferOut_long(2658) <= dataBufferIn_long(  78);
	dataBufferOut_long(3401) <= dataBufferIn_long(  79);
	dataBufferOut_long(4144) <= dataBufferIn_long(  80);
	dataBufferOut_long(4887) <= dataBufferIn_long(  81);
	dataBufferOut_long(5630) <= dataBufferIn_long(  82);
	dataBufferOut_long( 229) <= dataBufferIn_long(  83);
	dataBufferOut_long( 972) <= dataBufferIn_long(  84);
	dataBufferOut_long(1715) <= dataBufferIn_long(  85);
	dataBufferOut_long(2458) <= dataBufferIn_long(  86);
	dataBufferOut_long(3201) <= dataBufferIn_long(  87);
	dataBufferOut_long(3944) <= dataBufferIn_long(  88);
	dataBufferOut_long(4687) <= dataBufferIn_long(  89);
	dataBufferOut_long(5430) <= dataBufferIn_long(  90);
	dataBufferOut_long(  29) <= dataBufferIn_long(  91);
	dataBufferOut_long( 772) <= dataBufferIn_long(  92);
	dataBufferOut_long(1515) <= dataBufferIn_long(  93);
	dataBufferOut_long(2258) <= dataBufferIn_long(  94);
	dataBufferOut_long(3001) <= dataBufferIn_long(  95);
	dataBufferOut_long(3744) <= dataBufferIn_long(  96);
	dataBufferOut_long(4487) <= dataBufferIn_long(  97);
	dataBufferOut_long(5230) <= dataBufferIn_long(  98);
	dataBufferOut_long(5973) <= dataBufferIn_long(  99);
	dataBufferOut_long( 572) <= dataBufferIn_long( 100);
	dataBufferOut_long(1315) <= dataBufferIn_long( 101);
	dataBufferOut_long(2058) <= dataBufferIn_long( 102);
	dataBufferOut_long(2801) <= dataBufferIn_long( 103);
	dataBufferOut_long(3544) <= dataBufferIn_long( 104);
	dataBufferOut_long(4287) <= dataBufferIn_long( 105);
	dataBufferOut_long(5030) <= dataBufferIn_long( 106);
	dataBufferOut_long(5773) <= dataBufferIn_long( 107);
	dataBufferOut_long( 372) <= dataBufferIn_long( 108);
	dataBufferOut_long(1115) <= dataBufferIn_long( 109);
	dataBufferOut_long(1858) <= dataBufferIn_long( 110);
	dataBufferOut_long(2601) <= dataBufferIn_long( 111);
	dataBufferOut_long(3344) <= dataBufferIn_long( 112);
	dataBufferOut_long(4087) <= dataBufferIn_long( 113);
	dataBufferOut_long(4830) <= dataBufferIn_long( 114);
	dataBufferOut_long(5573) <= dataBufferIn_long( 115);
	dataBufferOut_long( 172) <= dataBufferIn_long( 116);
	dataBufferOut_long( 915) <= dataBufferIn_long( 117);
	dataBufferOut_long(1658) <= dataBufferIn_long( 118);
	dataBufferOut_long(2401) <= dataBufferIn_long( 119);
	dataBufferOut_long(3144) <= dataBufferIn_long( 120);
	dataBufferOut_long(3887) <= dataBufferIn_long( 121);
	dataBufferOut_long(4630) <= dataBufferIn_long( 122);
	dataBufferOut_long(5373) <= dataBufferIn_long( 123);
	dataBufferOut_long(6116) <= dataBufferIn_long( 124);
	dataBufferOut_long( 715) <= dataBufferIn_long( 125);
	dataBufferOut_long(1458) <= dataBufferIn_long( 126);
	dataBufferOut_long(2201) <= dataBufferIn_long( 127);
	dataBufferOut_long(2944) <= dataBufferIn_long( 128);
	dataBufferOut_long(3687) <= dataBufferIn_long( 129);
	dataBufferOut_long(4430) <= dataBufferIn_long( 130);
	dataBufferOut_long(5173) <= dataBufferIn_long( 131);
	dataBufferOut_long(5916) <= dataBufferIn_long( 132);
	dataBufferOut_long( 515) <= dataBufferIn_long( 133);
	dataBufferOut_long(1258) <= dataBufferIn_long( 134);
	dataBufferOut_long(2001) <= dataBufferIn_long( 135);
	dataBufferOut_long(2744) <= dataBufferIn_long( 136);
	dataBufferOut_long(3487) <= dataBufferIn_long( 137);
	dataBufferOut_long(4230) <= dataBufferIn_long( 138);
	dataBufferOut_long(4973) <= dataBufferIn_long( 139);
	dataBufferOut_long(5716) <= dataBufferIn_long( 140);
	dataBufferOut_long( 315) <= dataBufferIn_long( 141);
	dataBufferOut_long(1058) <= dataBufferIn_long( 142);
	dataBufferOut_long(1801) <= dataBufferIn_long( 143);
	dataBufferOut_long(2544) <= dataBufferIn_long( 144);
	dataBufferOut_long(3287) <= dataBufferIn_long( 145);
	dataBufferOut_long(4030) <= dataBufferIn_long( 146);
	dataBufferOut_long(4773) <= dataBufferIn_long( 147);
	dataBufferOut_long(5516) <= dataBufferIn_long( 148);
	dataBufferOut_long( 115) <= dataBufferIn_long( 149);
	dataBufferOut_long( 858) <= dataBufferIn_long( 150);
	dataBufferOut_long(1601) <= dataBufferIn_long( 151);
	dataBufferOut_long(2344) <= dataBufferIn_long( 152);
	dataBufferOut_long(3087) <= dataBufferIn_long( 153);
	dataBufferOut_long(3830) <= dataBufferIn_long( 154);
	dataBufferOut_long(4573) <= dataBufferIn_long( 155);
	dataBufferOut_long(5316) <= dataBufferIn_long( 156);
	dataBufferOut_long(6059) <= dataBufferIn_long( 157);
	dataBufferOut_long( 658) <= dataBufferIn_long( 158);
	dataBufferOut_long(1401) <= dataBufferIn_long( 159);
	dataBufferOut_long(2144) <= dataBufferIn_long( 160);
	dataBufferOut_long(2887) <= dataBufferIn_long( 161);
	dataBufferOut_long(3630) <= dataBufferIn_long( 162);
	dataBufferOut_long(4373) <= dataBufferIn_long( 163);
	dataBufferOut_long(5116) <= dataBufferIn_long( 164);
	dataBufferOut_long(5859) <= dataBufferIn_long( 165);
	dataBufferOut_long( 458) <= dataBufferIn_long( 166);
	dataBufferOut_long(1201) <= dataBufferIn_long( 167);
	dataBufferOut_long(1944) <= dataBufferIn_long( 168);
	dataBufferOut_long(2687) <= dataBufferIn_long( 169);
	dataBufferOut_long(3430) <= dataBufferIn_long( 170);
	dataBufferOut_long(4173) <= dataBufferIn_long( 171);
	dataBufferOut_long(4916) <= dataBufferIn_long( 172);
	dataBufferOut_long(5659) <= dataBufferIn_long( 173);
	dataBufferOut_long( 258) <= dataBufferIn_long( 174);
	dataBufferOut_long(1001) <= dataBufferIn_long( 175);
	dataBufferOut_long(1744) <= dataBufferIn_long( 176);
	dataBufferOut_long(2487) <= dataBufferIn_long( 177);
	dataBufferOut_long(3230) <= dataBufferIn_long( 178);
	dataBufferOut_long(3973) <= dataBufferIn_long( 179);
	dataBufferOut_long(4716) <= dataBufferIn_long( 180);
	dataBufferOut_long(5459) <= dataBufferIn_long( 181);
	dataBufferOut_long(  58) <= dataBufferIn_long( 182);
	dataBufferOut_long( 801) <= dataBufferIn_long( 183);
	dataBufferOut_long(1544) <= dataBufferIn_long( 184);
	dataBufferOut_long(2287) <= dataBufferIn_long( 185);
	dataBufferOut_long(3030) <= dataBufferIn_long( 186);
	dataBufferOut_long(3773) <= dataBufferIn_long( 187);
	dataBufferOut_long(4516) <= dataBufferIn_long( 188);
	dataBufferOut_long(5259) <= dataBufferIn_long( 189);
	dataBufferOut_long(6002) <= dataBufferIn_long( 190);
	dataBufferOut_long( 601) <= dataBufferIn_long( 191);
	dataBufferOut_long(1344) <= dataBufferIn_long( 192);
	dataBufferOut_long(2087) <= dataBufferIn_long( 193);
	dataBufferOut_long(2830) <= dataBufferIn_long( 194);
	dataBufferOut_long(3573) <= dataBufferIn_long( 195);
	dataBufferOut_long(4316) <= dataBufferIn_long( 196);
	dataBufferOut_long(5059) <= dataBufferIn_long( 197);
	dataBufferOut_long(5802) <= dataBufferIn_long( 198);
	dataBufferOut_long( 401) <= dataBufferIn_long( 199);
	dataBufferOut_long(1144) <= dataBufferIn_long( 200);
	dataBufferOut_long(1887) <= dataBufferIn_long( 201);
	dataBufferOut_long(2630) <= dataBufferIn_long( 202);
	dataBufferOut_long(3373) <= dataBufferIn_long( 203);
	dataBufferOut_long(4116) <= dataBufferIn_long( 204);
	dataBufferOut_long(4859) <= dataBufferIn_long( 205);
	dataBufferOut_long(5602) <= dataBufferIn_long( 206);
	dataBufferOut_long( 201) <= dataBufferIn_long( 207);
	dataBufferOut_long( 944) <= dataBufferIn_long( 208);
	dataBufferOut_long(1687) <= dataBufferIn_long( 209);
	dataBufferOut_long(2430) <= dataBufferIn_long( 210);
	dataBufferOut_long(3173) <= dataBufferIn_long( 211);
	dataBufferOut_long(3916) <= dataBufferIn_long( 212);
	dataBufferOut_long(4659) <= dataBufferIn_long( 213);
	dataBufferOut_long(5402) <= dataBufferIn_long( 214);
	dataBufferOut_long(   1) <= dataBufferIn_long( 215);
	dataBufferOut_long( 744) <= dataBufferIn_long( 216);
	dataBufferOut_long(1487) <= dataBufferIn_long( 217);
	dataBufferOut_long(2230) <= dataBufferIn_long( 218);
	dataBufferOut_long(2973) <= dataBufferIn_long( 219);
	dataBufferOut_long(3716) <= dataBufferIn_long( 220);
	dataBufferOut_long(4459) <= dataBufferIn_long( 221);
	dataBufferOut_long(5202) <= dataBufferIn_long( 222);
	dataBufferOut_long(5945) <= dataBufferIn_long( 223);
	dataBufferOut_long( 544) <= dataBufferIn_long( 224);
	dataBufferOut_long(1287) <= dataBufferIn_long( 225);
	dataBufferOut_long(2030) <= dataBufferIn_long( 226);
	dataBufferOut_long(2773) <= dataBufferIn_long( 227);
	dataBufferOut_long(3516) <= dataBufferIn_long( 228);
	dataBufferOut_long(4259) <= dataBufferIn_long( 229);
	dataBufferOut_long(5002) <= dataBufferIn_long( 230);
	dataBufferOut_long(5745) <= dataBufferIn_long( 231);
	dataBufferOut_long( 344) <= dataBufferIn_long( 232);
	dataBufferOut_long(1087) <= dataBufferIn_long( 233);
	dataBufferOut_long(1830) <= dataBufferIn_long( 234);
	dataBufferOut_long(2573) <= dataBufferIn_long( 235);
	dataBufferOut_long(3316) <= dataBufferIn_long( 236);
	dataBufferOut_long(4059) <= dataBufferIn_long( 237);
	dataBufferOut_long(4802) <= dataBufferIn_long( 238);
	dataBufferOut_long(5545) <= dataBufferIn_long( 239);
	dataBufferOut_long( 144) <= dataBufferIn_long( 240);
	dataBufferOut_long( 887) <= dataBufferIn_long( 241);
	dataBufferOut_long(1630) <= dataBufferIn_long( 242);
	dataBufferOut_long(2373) <= dataBufferIn_long( 243);
	dataBufferOut_long(3116) <= dataBufferIn_long( 244);
	dataBufferOut_long(3859) <= dataBufferIn_long( 245);
	dataBufferOut_long(4602) <= dataBufferIn_long( 246);
	dataBufferOut_long(5345) <= dataBufferIn_long( 247);
	dataBufferOut_long(6088) <= dataBufferIn_long( 248);
	dataBufferOut_long( 687) <= dataBufferIn_long( 249);
	dataBufferOut_long(1430) <= dataBufferIn_long( 250);
	dataBufferOut_long(2173) <= dataBufferIn_long( 251);
	dataBufferOut_long(2916) <= dataBufferIn_long( 252);
	dataBufferOut_long(3659) <= dataBufferIn_long( 253);
	dataBufferOut_long(4402) <= dataBufferIn_long( 254);
	dataBufferOut_long(5145) <= dataBufferIn_long( 255);
	dataBufferOut_long(5888) <= dataBufferIn_long( 256);
	dataBufferOut_long( 487) <= dataBufferIn_long( 257);
	dataBufferOut_long(1230) <= dataBufferIn_long( 258);
	dataBufferOut_long(1973) <= dataBufferIn_long( 259);
	dataBufferOut_long(2716) <= dataBufferIn_long( 260);
	dataBufferOut_long(3459) <= dataBufferIn_long( 261);
	dataBufferOut_long(4202) <= dataBufferIn_long( 262);
	dataBufferOut_long(4945) <= dataBufferIn_long( 263);
	dataBufferOut_long(5688) <= dataBufferIn_long( 264);
	dataBufferOut_long( 287) <= dataBufferIn_long( 265);
	dataBufferOut_long(1030) <= dataBufferIn_long( 266);
	dataBufferOut_long(1773) <= dataBufferIn_long( 267);
	dataBufferOut_long(2516) <= dataBufferIn_long( 268);
	dataBufferOut_long(3259) <= dataBufferIn_long( 269);
	dataBufferOut_long(4002) <= dataBufferIn_long( 270);
	dataBufferOut_long(4745) <= dataBufferIn_long( 271);
	dataBufferOut_long(5488) <= dataBufferIn_long( 272);
	dataBufferOut_long(  87) <= dataBufferIn_long( 273);
	dataBufferOut_long( 830) <= dataBufferIn_long( 274);
	dataBufferOut_long(1573) <= dataBufferIn_long( 275);
	dataBufferOut_long(2316) <= dataBufferIn_long( 276);
	dataBufferOut_long(3059) <= dataBufferIn_long( 277);
	dataBufferOut_long(3802) <= dataBufferIn_long( 278);
	dataBufferOut_long(4545) <= dataBufferIn_long( 279);
	dataBufferOut_long(5288) <= dataBufferIn_long( 280);
	dataBufferOut_long(6031) <= dataBufferIn_long( 281);
	dataBufferOut_long( 630) <= dataBufferIn_long( 282);
	dataBufferOut_long(1373) <= dataBufferIn_long( 283);
	dataBufferOut_long(2116) <= dataBufferIn_long( 284);
	dataBufferOut_long(2859) <= dataBufferIn_long( 285);
	dataBufferOut_long(3602) <= dataBufferIn_long( 286);
	dataBufferOut_long(4345) <= dataBufferIn_long( 287);
	dataBufferOut_long(5088) <= dataBufferIn_long( 288);
	dataBufferOut_long(5831) <= dataBufferIn_long( 289);
	dataBufferOut_long( 430) <= dataBufferIn_long( 290);
	dataBufferOut_long(1173) <= dataBufferIn_long( 291);
	dataBufferOut_long(1916) <= dataBufferIn_long( 292);
	dataBufferOut_long(2659) <= dataBufferIn_long( 293);
	dataBufferOut_long(3402) <= dataBufferIn_long( 294);
	dataBufferOut_long(4145) <= dataBufferIn_long( 295);
	dataBufferOut_long(4888) <= dataBufferIn_long( 296);
	dataBufferOut_long(5631) <= dataBufferIn_long( 297);
	dataBufferOut_long( 230) <= dataBufferIn_long( 298);
	dataBufferOut_long( 973) <= dataBufferIn_long( 299);
	dataBufferOut_long(1716) <= dataBufferIn_long( 300);
	dataBufferOut_long(2459) <= dataBufferIn_long( 301);
	dataBufferOut_long(3202) <= dataBufferIn_long( 302);
	dataBufferOut_long(3945) <= dataBufferIn_long( 303);
	dataBufferOut_long(4688) <= dataBufferIn_long( 304);
	dataBufferOut_long(5431) <= dataBufferIn_long( 305);
	dataBufferOut_long(  30) <= dataBufferIn_long( 306);
	dataBufferOut_long( 773) <= dataBufferIn_long( 307);
	dataBufferOut_long(1516) <= dataBufferIn_long( 308);
	dataBufferOut_long(2259) <= dataBufferIn_long( 309);
	dataBufferOut_long(3002) <= dataBufferIn_long( 310);
	dataBufferOut_long(3745) <= dataBufferIn_long( 311);
	dataBufferOut_long(4488) <= dataBufferIn_long( 312);
	dataBufferOut_long(5231) <= dataBufferIn_long( 313);
	dataBufferOut_long(5974) <= dataBufferIn_long( 314);
	dataBufferOut_long( 573) <= dataBufferIn_long( 315);
	dataBufferOut_long(1316) <= dataBufferIn_long( 316);
	dataBufferOut_long(2059) <= dataBufferIn_long( 317);
	dataBufferOut_long(2802) <= dataBufferIn_long( 318);
	dataBufferOut_long(3545) <= dataBufferIn_long( 319);
	dataBufferOut_long(4288) <= dataBufferIn_long( 320);
	dataBufferOut_long(5031) <= dataBufferIn_long( 321);
	dataBufferOut_long(5774) <= dataBufferIn_long( 322);
	dataBufferOut_long( 373) <= dataBufferIn_long( 323);
	dataBufferOut_long(1116) <= dataBufferIn_long( 324);
	dataBufferOut_long(1859) <= dataBufferIn_long( 325);
	dataBufferOut_long(2602) <= dataBufferIn_long( 326);
	dataBufferOut_long(3345) <= dataBufferIn_long( 327);
	dataBufferOut_long(4088) <= dataBufferIn_long( 328);
	dataBufferOut_long(4831) <= dataBufferIn_long( 329);
	dataBufferOut_long(5574) <= dataBufferIn_long( 330);
	dataBufferOut_long( 173) <= dataBufferIn_long( 331);
	dataBufferOut_long( 916) <= dataBufferIn_long( 332);
	dataBufferOut_long(1659) <= dataBufferIn_long( 333);
	dataBufferOut_long(2402) <= dataBufferIn_long( 334);
	dataBufferOut_long(3145) <= dataBufferIn_long( 335);
	dataBufferOut_long(3888) <= dataBufferIn_long( 336);
	dataBufferOut_long(4631) <= dataBufferIn_long( 337);
	dataBufferOut_long(5374) <= dataBufferIn_long( 338);
	dataBufferOut_long(6117) <= dataBufferIn_long( 339);
	dataBufferOut_long( 716) <= dataBufferIn_long( 340);
	dataBufferOut_long(1459) <= dataBufferIn_long( 341);
	dataBufferOut_long(2202) <= dataBufferIn_long( 342);
	dataBufferOut_long(2945) <= dataBufferIn_long( 343);
	dataBufferOut_long(3688) <= dataBufferIn_long( 344);
	dataBufferOut_long(4431) <= dataBufferIn_long( 345);
	dataBufferOut_long(5174) <= dataBufferIn_long( 346);
	dataBufferOut_long(5917) <= dataBufferIn_long( 347);
	dataBufferOut_long( 516) <= dataBufferIn_long( 348);
	dataBufferOut_long(1259) <= dataBufferIn_long( 349);
	dataBufferOut_long(2002) <= dataBufferIn_long( 350);
	dataBufferOut_long(2745) <= dataBufferIn_long( 351);
	dataBufferOut_long(3488) <= dataBufferIn_long( 352);
	dataBufferOut_long(4231) <= dataBufferIn_long( 353);
	dataBufferOut_long(4974) <= dataBufferIn_long( 354);
	dataBufferOut_long(5717) <= dataBufferIn_long( 355);
	dataBufferOut_long( 316) <= dataBufferIn_long( 356);
	dataBufferOut_long(1059) <= dataBufferIn_long( 357);
	dataBufferOut_long(1802) <= dataBufferIn_long( 358);
	dataBufferOut_long(2545) <= dataBufferIn_long( 359);
	dataBufferOut_long(3288) <= dataBufferIn_long( 360);
	dataBufferOut_long(4031) <= dataBufferIn_long( 361);
	dataBufferOut_long(4774) <= dataBufferIn_long( 362);
	dataBufferOut_long(5517) <= dataBufferIn_long( 363);
	dataBufferOut_long( 116) <= dataBufferIn_long( 364);
	dataBufferOut_long( 859) <= dataBufferIn_long( 365);
	dataBufferOut_long(1602) <= dataBufferIn_long( 366);
	dataBufferOut_long(2345) <= dataBufferIn_long( 367);
	dataBufferOut_long(3088) <= dataBufferIn_long( 368);
	dataBufferOut_long(3831) <= dataBufferIn_long( 369);
	dataBufferOut_long(4574) <= dataBufferIn_long( 370);
	dataBufferOut_long(5317) <= dataBufferIn_long( 371);
	dataBufferOut_long(6060) <= dataBufferIn_long( 372);
	dataBufferOut_long( 659) <= dataBufferIn_long( 373);
	dataBufferOut_long(1402) <= dataBufferIn_long( 374);
	dataBufferOut_long(2145) <= dataBufferIn_long( 375);
	dataBufferOut_long(2888) <= dataBufferIn_long( 376);
	dataBufferOut_long(3631) <= dataBufferIn_long( 377);
	dataBufferOut_long(4374) <= dataBufferIn_long( 378);
	dataBufferOut_long(5117) <= dataBufferIn_long( 379);
	dataBufferOut_long(5860) <= dataBufferIn_long( 380);
	dataBufferOut_long( 459) <= dataBufferIn_long( 381);
	dataBufferOut_long(1202) <= dataBufferIn_long( 382);
	dataBufferOut_long(1945) <= dataBufferIn_long( 383);
	dataBufferOut_long(2688) <= dataBufferIn_long( 384);
	dataBufferOut_long(3431) <= dataBufferIn_long( 385);
	dataBufferOut_long(4174) <= dataBufferIn_long( 386);
	dataBufferOut_long(4917) <= dataBufferIn_long( 387);
	dataBufferOut_long(5660) <= dataBufferIn_long( 388);
	dataBufferOut_long( 259) <= dataBufferIn_long( 389);
	dataBufferOut_long(1002) <= dataBufferIn_long( 390);
	dataBufferOut_long(1745) <= dataBufferIn_long( 391);
	dataBufferOut_long(2488) <= dataBufferIn_long( 392);
	dataBufferOut_long(3231) <= dataBufferIn_long( 393);
	dataBufferOut_long(3974) <= dataBufferIn_long( 394);
	dataBufferOut_long(4717) <= dataBufferIn_long( 395);
	dataBufferOut_long(5460) <= dataBufferIn_long( 396);
	dataBufferOut_long(  59) <= dataBufferIn_long( 397);
	dataBufferOut_long( 802) <= dataBufferIn_long( 398);
	dataBufferOut_long(1545) <= dataBufferIn_long( 399);
	dataBufferOut_long(2288) <= dataBufferIn_long( 400);
	dataBufferOut_long(3031) <= dataBufferIn_long( 401);
	dataBufferOut_long(3774) <= dataBufferIn_long( 402);
	dataBufferOut_long(4517) <= dataBufferIn_long( 403);
	dataBufferOut_long(5260) <= dataBufferIn_long( 404);
	dataBufferOut_long(6003) <= dataBufferIn_long( 405);
	dataBufferOut_long( 602) <= dataBufferIn_long( 406);
	dataBufferOut_long(1345) <= dataBufferIn_long( 407);
	dataBufferOut_long(2088) <= dataBufferIn_long( 408);
	dataBufferOut_long(2831) <= dataBufferIn_long( 409);
	dataBufferOut_long(3574) <= dataBufferIn_long( 410);
	dataBufferOut_long(4317) <= dataBufferIn_long( 411);
	dataBufferOut_long(5060) <= dataBufferIn_long( 412);
	dataBufferOut_long(5803) <= dataBufferIn_long( 413);
	dataBufferOut_long( 402) <= dataBufferIn_long( 414);
	dataBufferOut_long(1145) <= dataBufferIn_long( 415);
	dataBufferOut_long(1888) <= dataBufferIn_long( 416);
	dataBufferOut_long(2631) <= dataBufferIn_long( 417);
	dataBufferOut_long(3374) <= dataBufferIn_long( 418);
	dataBufferOut_long(4117) <= dataBufferIn_long( 419);
	dataBufferOut_long(4860) <= dataBufferIn_long( 420);
	dataBufferOut_long(5603) <= dataBufferIn_long( 421);
	dataBufferOut_long( 202) <= dataBufferIn_long( 422);
	dataBufferOut_long( 945) <= dataBufferIn_long( 423);
	dataBufferOut_long(1688) <= dataBufferIn_long( 424);
	dataBufferOut_long(2431) <= dataBufferIn_long( 425);
	dataBufferOut_long(3174) <= dataBufferIn_long( 426);
	dataBufferOut_long(3917) <= dataBufferIn_long( 427);
	dataBufferOut_long(4660) <= dataBufferIn_long( 428);
	dataBufferOut_long(5403) <= dataBufferIn_long( 429);
	dataBufferOut_long(   2) <= dataBufferIn_long( 430);
	dataBufferOut_long( 745) <= dataBufferIn_long( 431);
	dataBufferOut_long(1488) <= dataBufferIn_long( 432);
	dataBufferOut_long(2231) <= dataBufferIn_long( 433);
	dataBufferOut_long(2974) <= dataBufferIn_long( 434);
	dataBufferOut_long(3717) <= dataBufferIn_long( 435);
	dataBufferOut_long(4460) <= dataBufferIn_long( 436);
	dataBufferOut_long(5203) <= dataBufferIn_long( 437);
	dataBufferOut_long(5946) <= dataBufferIn_long( 438);
	dataBufferOut_long( 545) <= dataBufferIn_long( 439);
	dataBufferOut_long(1288) <= dataBufferIn_long( 440);
	dataBufferOut_long(2031) <= dataBufferIn_long( 441);
	dataBufferOut_long(2774) <= dataBufferIn_long( 442);
	dataBufferOut_long(3517) <= dataBufferIn_long( 443);
	dataBufferOut_long(4260) <= dataBufferIn_long( 444);
	dataBufferOut_long(5003) <= dataBufferIn_long( 445);
	dataBufferOut_long(5746) <= dataBufferIn_long( 446);
	dataBufferOut_long( 345) <= dataBufferIn_long( 447);
	dataBufferOut_long(1088) <= dataBufferIn_long( 448);
	dataBufferOut_long(1831) <= dataBufferIn_long( 449);
	dataBufferOut_long(2574) <= dataBufferIn_long( 450);
	dataBufferOut_long(3317) <= dataBufferIn_long( 451);
	dataBufferOut_long(4060) <= dataBufferIn_long( 452);
	dataBufferOut_long(4803) <= dataBufferIn_long( 453);
	dataBufferOut_long(5546) <= dataBufferIn_long( 454);
	dataBufferOut_long( 145) <= dataBufferIn_long( 455);
	dataBufferOut_long( 888) <= dataBufferIn_long( 456);
	dataBufferOut_long(1631) <= dataBufferIn_long( 457);
	dataBufferOut_long(2374) <= dataBufferIn_long( 458);
	dataBufferOut_long(3117) <= dataBufferIn_long( 459);
	dataBufferOut_long(3860) <= dataBufferIn_long( 460);
	dataBufferOut_long(4603) <= dataBufferIn_long( 461);
	dataBufferOut_long(5346) <= dataBufferIn_long( 462);
	dataBufferOut_long(6089) <= dataBufferIn_long( 463);
	dataBufferOut_long( 688) <= dataBufferIn_long( 464);
	dataBufferOut_long(1431) <= dataBufferIn_long( 465);
	dataBufferOut_long(2174) <= dataBufferIn_long( 466);
	dataBufferOut_long(2917) <= dataBufferIn_long( 467);
	dataBufferOut_long(3660) <= dataBufferIn_long( 468);
	dataBufferOut_long(4403) <= dataBufferIn_long( 469);
	dataBufferOut_long(5146) <= dataBufferIn_long( 470);
	dataBufferOut_long(5889) <= dataBufferIn_long( 471);
	dataBufferOut_long( 488) <= dataBufferIn_long( 472);
	dataBufferOut_long(1231) <= dataBufferIn_long( 473);
	dataBufferOut_long(1974) <= dataBufferIn_long( 474);
	dataBufferOut_long(2717) <= dataBufferIn_long( 475);
	dataBufferOut_long(3460) <= dataBufferIn_long( 476);
	dataBufferOut_long(4203) <= dataBufferIn_long( 477);
	dataBufferOut_long(4946) <= dataBufferIn_long( 478);
	dataBufferOut_long(5689) <= dataBufferIn_long( 479);
	dataBufferOut_long( 288) <= dataBufferIn_long( 480);
	dataBufferOut_long(1031) <= dataBufferIn_long( 481);
	dataBufferOut_long(1774) <= dataBufferIn_long( 482);
	dataBufferOut_long(2517) <= dataBufferIn_long( 483);
	dataBufferOut_long(3260) <= dataBufferIn_long( 484);
	dataBufferOut_long(4003) <= dataBufferIn_long( 485);
	dataBufferOut_long(4746) <= dataBufferIn_long( 486);
	dataBufferOut_long(5489) <= dataBufferIn_long( 487);
	dataBufferOut_long(  88) <= dataBufferIn_long( 488);
	dataBufferOut_long( 831) <= dataBufferIn_long( 489);
	dataBufferOut_long(1574) <= dataBufferIn_long( 490);
	dataBufferOut_long(2317) <= dataBufferIn_long( 491);
	dataBufferOut_long(3060) <= dataBufferIn_long( 492);
	dataBufferOut_long(3803) <= dataBufferIn_long( 493);
	dataBufferOut_long(4546) <= dataBufferIn_long( 494);
	dataBufferOut_long(5289) <= dataBufferIn_long( 495);
	dataBufferOut_long(6032) <= dataBufferIn_long( 496);
	dataBufferOut_long( 631) <= dataBufferIn_long( 497);
	dataBufferOut_long(1374) <= dataBufferIn_long( 498);
	dataBufferOut_long(2117) <= dataBufferIn_long( 499);
	dataBufferOut_long(2860) <= dataBufferIn_long( 500);
	dataBufferOut_long(3603) <= dataBufferIn_long( 501);
	dataBufferOut_long(4346) <= dataBufferIn_long( 502);
	dataBufferOut_long(5089) <= dataBufferIn_long( 503);
	dataBufferOut_long(5832) <= dataBufferIn_long( 504);
	dataBufferOut_long( 431) <= dataBufferIn_long( 505);
	dataBufferOut_long(1174) <= dataBufferIn_long( 506);
	dataBufferOut_long(1917) <= dataBufferIn_long( 507);
	dataBufferOut_long(2660) <= dataBufferIn_long( 508);
	dataBufferOut_long(3403) <= dataBufferIn_long( 509);
	dataBufferOut_long(4146) <= dataBufferIn_long( 510);
	dataBufferOut_long(4889) <= dataBufferIn_long( 511);
	dataBufferOut_long(5632) <= dataBufferIn_long( 512);
	dataBufferOut_long( 231) <= dataBufferIn_long( 513);
	dataBufferOut_long( 974) <= dataBufferIn_long( 514);
	dataBufferOut_long(1717) <= dataBufferIn_long( 515);
	dataBufferOut_long(2460) <= dataBufferIn_long( 516);
	dataBufferOut_long(3203) <= dataBufferIn_long( 517);
	dataBufferOut_long(3946) <= dataBufferIn_long( 518);
	dataBufferOut_long(4689) <= dataBufferIn_long( 519);
	dataBufferOut_long(5432) <= dataBufferIn_long( 520);
	dataBufferOut_long(  31) <= dataBufferIn_long( 521);
	dataBufferOut_long( 774) <= dataBufferIn_long( 522);
	dataBufferOut_long(1517) <= dataBufferIn_long( 523);
	dataBufferOut_long(2260) <= dataBufferIn_long( 524);
	dataBufferOut_long(3003) <= dataBufferIn_long( 525);
	dataBufferOut_long(3746) <= dataBufferIn_long( 526);
	dataBufferOut_long(4489) <= dataBufferIn_long( 527);
	dataBufferOut_long(5232) <= dataBufferIn_long( 528);
	dataBufferOut_long(5975) <= dataBufferIn_long( 529);
	dataBufferOut_long( 574) <= dataBufferIn_long( 530);
	dataBufferOut_long(1317) <= dataBufferIn_long( 531);
	dataBufferOut_long(2060) <= dataBufferIn_long( 532);
	dataBufferOut_long(2803) <= dataBufferIn_long( 533);
	dataBufferOut_long(3546) <= dataBufferIn_long( 534);
	dataBufferOut_long(4289) <= dataBufferIn_long( 535);
	dataBufferOut_long(5032) <= dataBufferIn_long( 536);
	dataBufferOut_long(5775) <= dataBufferIn_long( 537);
	dataBufferOut_long( 374) <= dataBufferIn_long( 538);
	dataBufferOut_long(1117) <= dataBufferIn_long( 539);
	dataBufferOut_long(1860) <= dataBufferIn_long( 540);
	dataBufferOut_long(2603) <= dataBufferIn_long( 541);
	dataBufferOut_long(3346) <= dataBufferIn_long( 542);
	dataBufferOut_long(4089) <= dataBufferIn_long( 543);
	dataBufferOut_long(4832) <= dataBufferIn_long( 544);
	dataBufferOut_long(5575) <= dataBufferIn_long( 545);
	dataBufferOut_long( 174) <= dataBufferIn_long( 546);
	dataBufferOut_long( 917) <= dataBufferIn_long( 547);
	dataBufferOut_long(1660) <= dataBufferIn_long( 548);
	dataBufferOut_long(2403) <= dataBufferIn_long( 549);
	dataBufferOut_long(3146) <= dataBufferIn_long( 550);
	dataBufferOut_long(3889) <= dataBufferIn_long( 551);
	dataBufferOut_long(4632) <= dataBufferIn_long( 552);
	dataBufferOut_long(5375) <= dataBufferIn_long( 553);
	dataBufferOut_long(6118) <= dataBufferIn_long( 554);
	dataBufferOut_long( 717) <= dataBufferIn_long( 555);
	dataBufferOut_long(1460) <= dataBufferIn_long( 556);
	dataBufferOut_long(2203) <= dataBufferIn_long( 557);
	dataBufferOut_long(2946) <= dataBufferIn_long( 558);
	dataBufferOut_long(3689) <= dataBufferIn_long( 559);
	dataBufferOut_long(4432) <= dataBufferIn_long( 560);
	dataBufferOut_long(5175) <= dataBufferIn_long( 561);
	dataBufferOut_long(5918) <= dataBufferIn_long( 562);
	dataBufferOut_long( 517) <= dataBufferIn_long( 563);
	dataBufferOut_long(1260) <= dataBufferIn_long( 564);
	dataBufferOut_long(2003) <= dataBufferIn_long( 565);
	dataBufferOut_long(2746) <= dataBufferIn_long( 566);
	dataBufferOut_long(3489) <= dataBufferIn_long( 567);
	dataBufferOut_long(4232) <= dataBufferIn_long( 568);
	dataBufferOut_long(4975) <= dataBufferIn_long( 569);
	dataBufferOut_long(5718) <= dataBufferIn_long( 570);
	dataBufferOut_long( 317) <= dataBufferIn_long( 571);
	dataBufferOut_long(1060) <= dataBufferIn_long( 572);
	dataBufferOut_long(1803) <= dataBufferIn_long( 573);
	dataBufferOut_long(2546) <= dataBufferIn_long( 574);
	dataBufferOut_long(3289) <= dataBufferIn_long( 575);
	dataBufferOut_long(4032) <= dataBufferIn_long( 576);
	dataBufferOut_long(4775) <= dataBufferIn_long( 577);
	dataBufferOut_long(5518) <= dataBufferIn_long( 578);
	dataBufferOut_long( 117) <= dataBufferIn_long( 579);
	dataBufferOut_long( 860) <= dataBufferIn_long( 580);
	dataBufferOut_long(1603) <= dataBufferIn_long( 581);
	dataBufferOut_long(2346) <= dataBufferIn_long( 582);
	dataBufferOut_long(3089) <= dataBufferIn_long( 583);
	dataBufferOut_long(3832) <= dataBufferIn_long( 584);
	dataBufferOut_long(4575) <= dataBufferIn_long( 585);
	dataBufferOut_long(5318) <= dataBufferIn_long( 586);
	dataBufferOut_long(6061) <= dataBufferIn_long( 587);
	dataBufferOut_long( 660) <= dataBufferIn_long( 588);
	dataBufferOut_long(1403) <= dataBufferIn_long( 589);
	dataBufferOut_long(2146) <= dataBufferIn_long( 590);
	dataBufferOut_long(2889) <= dataBufferIn_long( 591);
	dataBufferOut_long(3632) <= dataBufferIn_long( 592);
	dataBufferOut_long(4375) <= dataBufferIn_long( 593);
	dataBufferOut_long(5118) <= dataBufferIn_long( 594);
	dataBufferOut_long(5861) <= dataBufferIn_long( 595);
	dataBufferOut_long( 460) <= dataBufferIn_long( 596);
	dataBufferOut_long(1203) <= dataBufferIn_long( 597);
	dataBufferOut_long(1946) <= dataBufferIn_long( 598);
	dataBufferOut_long(2689) <= dataBufferIn_long( 599);
	dataBufferOut_long(3432) <= dataBufferIn_long( 600);
	dataBufferOut_long(4175) <= dataBufferIn_long( 601);
	dataBufferOut_long(4918) <= dataBufferIn_long( 602);
	dataBufferOut_long(5661) <= dataBufferIn_long( 603);
	dataBufferOut_long( 260) <= dataBufferIn_long( 604);
	dataBufferOut_long(1003) <= dataBufferIn_long( 605);
	dataBufferOut_long(1746) <= dataBufferIn_long( 606);
	dataBufferOut_long(2489) <= dataBufferIn_long( 607);
	dataBufferOut_long(3232) <= dataBufferIn_long( 608);
	dataBufferOut_long(3975) <= dataBufferIn_long( 609);
	dataBufferOut_long(4718) <= dataBufferIn_long( 610);
	dataBufferOut_long(5461) <= dataBufferIn_long( 611);
	dataBufferOut_long(  60) <= dataBufferIn_long( 612);
	dataBufferOut_long( 803) <= dataBufferIn_long( 613);
	dataBufferOut_long(1546) <= dataBufferIn_long( 614);
	dataBufferOut_long(2289) <= dataBufferIn_long( 615);
	dataBufferOut_long(3032) <= dataBufferIn_long( 616);
	dataBufferOut_long(3775) <= dataBufferIn_long( 617);
	dataBufferOut_long(4518) <= dataBufferIn_long( 618);
	dataBufferOut_long(5261) <= dataBufferIn_long( 619);
	dataBufferOut_long(6004) <= dataBufferIn_long( 620);
	dataBufferOut_long( 603) <= dataBufferIn_long( 621);
	dataBufferOut_long(1346) <= dataBufferIn_long( 622);
	dataBufferOut_long(2089) <= dataBufferIn_long( 623);
	dataBufferOut_long(2832) <= dataBufferIn_long( 624);
	dataBufferOut_long(3575) <= dataBufferIn_long( 625);
	dataBufferOut_long(4318) <= dataBufferIn_long( 626);
	dataBufferOut_long(5061) <= dataBufferIn_long( 627);
	dataBufferOut_long(5804) <= dataBufferIn_long( 628);
	dataBufferOut_long( 403) <= dataBufferIn_long( 629);
	dataBufferOut_long(1146) <= dataBufferIn_long( 630);
	dataBufferOut_long(1889) <= dataBufferIn_long( 631);
	dataBufferOut_long(2632) <= dataBufferIn_long( 632);
	dataBufferOut_long(3375) <= dataBufferIn_long( 633);
	dataBufferOut_long(4118) <= dataBufferIn_long( 634);
	dataBufferOut_long(4861) <= dataBufferIn_long( 635);
	dataBufferOut_long(5604) <= dataBufferIn_long( 636);
	dataBufferOut_long( 203) <= dataBufferIn_long( 637);
	dataBufferOut_long( 946) <= dataBufferIn_long( 638);
	dataBufferOut_long(1689) <= dataBufferIn_long( 639);
	dataBufferOut_long(2432) <= dataBufferIn_long( 640);
	dataBufferOut_long(3175) <= dataBufferIn_long( 641);
	dataBufferOut_long(3918) <= dataBufferIn_long( 642);
	dataBufferOut_long(4661) <= dataBufferIn_long( 643);
	dataBufferOut_long(5404) <= dataBufferIn_long( 644);
	dataBufferOut_long(   3) <= dataBufferIn_long( 645);
	dataBufferOut_long( 746) <= dataBufferIn_long( 646);
	dataBufferOut_long(1489) <= dataBufferIn_long( 647);
	dataBufferOut_long(2232) <= dataBufferIn_long( 648);
	dataBufferOut_long(2975) <= dataBufferIn_long( 649);
	dataBufferOut_long(3718) <= dataBufferIn_long( 650);
	dataBufferOut_long(4461) <= dataBufferIn_long( 651);
	dataBufferOut_long(5204) <= dataBufferIn_long( 652);
	dataBufferOut_long(5947) <= dataBufferIn_long( 653);
	dataBufferOut_long( 546) <= dataBufferIn_long( 654);
	dataBufferOut_long(1289) <= dataBufferIn_long( 655);
	dataBufferOut_long(2032) <= dataBufferIn_long( 656);
	dataBufferOut_long(2775) <= dataBufferIn_long( 657);
	dataBufferOut_long(3518) <= dataBufferIn_long( 658);
	dataBufferOut_long(4261) <= dataBufferIn_long( 659);
	dataBufferOut_long(5004) <= dataBufferIn_long( 660);
	dataBufferOut_long(5747) <= dataBufferIn_long( 661);
	dataBufferOut_long( 346) <= dataBufferIn_long( 662);
	dataBufferOut_long(1089) <= dataBufferIn_long( 663);
	dataBufferOut_long(1832) <= dataBufferIn_long( 664);
	dataBufferOut_long(2575) <= dataBufferIn_long( 665);
	dataBufferOut_long(3318) <= dataBufferIn_long( 666);
	dataBufferOut_long(4061) <= dataBufferIn_long( 667);
	dataBufferOut_long(4804) <= dataBufferIn_long( 668);
	dataBufferOut_long(5547) <= dataBufferIn_long( 669);
	dataBufferOut_long( 146) <= dataBufferIn_long( 670);
	dataBufferOut_long( 889) <= dataBufferIn_long( 671);
	dataBufferOut_long(1632) <= dataBufferIn_long( 672);
	dataBufferOut_long(2375) <= dataBufferIn_long( 673);
	dataBufferOut_long(3118) <= dataBufferIn_long( 674);
	dataBufferOut_long(3861) <= dataBufferIn_long( 675);
	dataBufferOut_long(4604) <= dataBufferIn_long( 676);
	dataBufferOut_long(5347) <= dataBufferIn_long( 677);
	dataBufferOut_long(6090) <= dataBufferIn_long( 678);
	dataBufferOut_long( 689) <= dataBufferIn_long( 679);
	dataBufferOut_long(1432) <= dataBufferIn_long( 680);
	dataBufferOut_long(2175) <= dataBufferIn_long( 681);
	dataBufferOut_long(2918) <= dataBufferIn_long( 682);
	dataBufferOut_long(3661) <= dataBufferIn_long( 683);
	dataBufferOut_long(4404) <= dataBufferIn_long( 684);
	dataBufferOut_long(5147) <= dataBufferIn_long( 685);
	dataBufferOut_long(5890) <= dataBufferIn_long( 686);
	dataBufferOut_long( 489) <= dataBufferIn_long( 687);
	dataBufferOut_long(1232) <= dataBufferIn_long( 688);
	dataBufferOut_long(1975) <= dataBufferIn_long( 689);
	dataBufferOut_long(2718) <= dataBufferIn_long( 690);
	dataBufferOut_long(3461) <= dataBufferIn_long( 691);
	dataBufferOut_long(4204) <= dataBufferIn_long( 692);
	dataBufferOut_long(4947) <= dataBufferIn_long( 693);
	dataBufferOut_long(5690) <= dataBufferIn_long( 694);
	dataBufferOut_long( 289) <= dataBufferIn_long( 695);
	dataBufferOut_long(1032) <= dataBufferIn_long( 696);
	dataBufferOut_long(1775) <= dataBufferIn_long( 697);
	dataBufferOut_long(2518) <= dataBufferIn_long( 698);
	dataBufferOut_long(3261) <= dataBufferIn_long( 699);
	dataBufferOut_long(4004) <= dataBufferIn_long( 700);
	dataBufferOut_long(4747) <= dataBufferIn_long( 701);
	dataBufferOut_long(5490) <= dataBufferIn_long( 702);
	dataBufferOut_long(  89) <= dataBufferIn_long( 703);
	dataBufferOut_long( 832) <= dataBufferIn_long( 704);
	dataBufferOut_long(1575) <= dataBufferIn_long( 705);
	dataBufferOut_long(2318) <= dataBufferIn_long( 706);
	dataBufferOut_long(3061) <= dataBufferIn_long( 707);
	dataBufferOut_long(3804) <= dataBufferIn_long( 708);
	dataBufferOut_long(4547) <= dataBufferIn_long( 709);
	dataBufferOut_long(5290) <= dataBufferIn_long( 710);
	dataBufferOut_long(6033) <= dataBufferIn_long( 711);
	dataBufferOut_long( 632) <= dataBufferIn_long( 712);
	dataBufferOut_long(1375) <= dataBufferIn_long( 713);
	dataBufferOut_long(2118) <= dataBufferIn_long( 714);
	dataBufferOut_long(2861) <= dataBufferIn_long( 715);
	dataBufferOut_long(3604) <= dataBufferIn_long( 716);
	dataBufferOut_long(4347) <= dataBufferIn_long( 717);
	dataBufferOut_long(5090) <= dataBufferIn_long( 718);
	dataBufferOut_long(5833) <= dataBufferIn_long( 719);
	dataBufferOut_long( 432) <= dataBufferIn_long( 720);
	dataBufferOut_long(1175) <= dataBufferIn_long( 721);
	dataBufferOut_long(1918) <= dataBufferIn_long( 722);
	dataBufferOut_long(2661) <= dataBufferIn_long( 723);
	dataBufferOut_long(3404) <= dataBufferIn_long( 724);
	dataBufferOut_long(4147) <= dataBufferIn_long( 725);
	dataBufferOut_long(4890) <= dataBufferIn_long( 726);
	dataBufferOut_long(5633) <= dataBufferIn_long( 727);
	dataBufferOut_long( 232) <= dataBufferIn_long( 728);
	dataBufferOut_long( 975) <= dataBufferIn_long( 729);
	dataBufferOut_long(1718) <= dataBufferIn_long( 730);
	dataBufferOut_long(2461) <= dataBufferIn_long( 731);
	dataBufferOut_long(3204) <= dataBufferIn_long( 732);
	dataBufferOut_long(3947) <= dataBufferIn_long( 733);
	dataBufferOut_long(4690) <= dataBufferIn_long( 734);
	dataBufferOut_long(5433) <= dataBufferIn_long( 735);
	dataBufferOut_long(  32) <= dataBufferIn_long( 736);
	dataBufferOut_long( 775) <= dataBufferIn_long( 737);
	dataBufferOut_long(1518) <= dataBufferIn_long( 738);
	dataBufferOut_long(2261) <= dataBufferIn_long( 739);
	dataBufferOut_long(3004) <= dataBufferIn_long( 740);
	dataBufferOut_long(3747) <= dataBufferIn_long( 741);
	dataBufferOut_long(4490) <= dataBufferIn_long( 742);
	dataBufferOut_long(5233) <= dataBufferIn_long( 743);
	dataBufferOut_long(5976) <= dataBufferIn_long( 744);
	dataBufferOut_long( 575) <= dataBufferIn_long( 745);
	dataBufferOut_long(1318) <= dataBufferIn_long( 746);
	dataBufferOut_long(2061) <= dataBufferIn_long( 747);
	dataBufferOut_long(2804) <= dataBufferIn_long( 748);
	dataBufferOut_long(3547) <= dataBufferIn_long( 749);
	dataBufferOut_long(4290) <= dataBufferIn_long( 750);
	dataBufferOut_long(5033) <= dataBufferIn_long( 751);
	dataBufferOut_long(5776) <= dataBufferIn_long( 752);
	dataBufferOut_long( 375) <= dataBufferIn_long( 753);
	dataBufferOut_long(1118) <= dataBufferIn_long( 754);
	dataBufferOut_long(1861) <= dataBufferIn_long( 755);
	dataBufferOut_long(2604) <= dataBufferIn_long( 756);
	dataBufferOut_long(3347) <= dataBufferIn_long( 757);
	dataBufferOut_long(4090) <= dataBufferIn_long( 758);
	dataBufferOut_long(4833) <= dataBufferIn_long( 759);
	dataBufferOut_long(5576) <= dataBufferIn_long( 760);
	dataBufferOut_long( 175) <= dataBufferIn_long( 761);
	dataBufferOut_long( 918) <= dataBufferIn_long( 762);
	dataBufferOut_long(1661) <= dataBufferIn_long( 763);
	dataBufferOut_long(2404) <= dataBufferIn_long( 764);
	dataBufferOut_long(3147) <= dataBufferIn_long( 765);
	dataBufferOut_long(3890) <= dataBufferIn_long( 766);
	dataBufferOut_long(4633) <= dataBufferIn_long( 767);
	dataBufferOut_long(5376) <= dataBufferIn_long( 768);
	dataBufferOut_long(6119) <= dataBufferIn_long( 769);
	dataBufferOut_long( 718) <= dataBufferIn_long( 770);
	dataBufferOut_long(1461) <= dataBufferIn_long( 771);
	dataBufferOut_long(2204) <= dataBufferIn_long( 772);
	dataBufferOut_long(2947) <= dataBufferIn_long( 773);
	dataBufferOut_long(3690) <= dataBufferIn_long( 774);
	dataBufferOut_long(4433) <= dataBufferIn_long( 775);
	dataBufferOut_long(5176) <= dataBufferIn_long( 776);
	dataBufferOut_long(5919) <= dataBufferIn_long( 777);
	dataBufferOut_long( 518) <= dataBufferIn_long( 778);
	dataBufferOut_long(1261) <= dataBufferIn_long( 779);
	dataBufferOut_long(2004) <= dataBufferIn_long( 780);
	dataBufferOut_long(2747) <= dataBufferIn_long( 781);
	dataBufferOut_long(3490) <= dataBufferIn_long( 782);
	dataBufferOut_long(4233) <= dataBufferIn_long( 783);
	dataBufferOut_long(4976) <= dataBufferIn_long( 784);
	dataBufferOut_long(5719) <= dataBufferIn_long( 785);
	dataBufferOut_long( 318) <= dataBufferIn_long( 786);
	dataBufferOut_long(1061) <= dataBufferIn_long( 787);
	dataBufferOut_long(1804) <= dataBufferIn_long( 788);
	dataBufferOut_long(2547) <= dataBufferIn_long( 789);
	dataBufferOut_long(3290) <= dataBufferIn_long( 790);
	dataBufferOut_long(4033) <= dataBufferIn_long( 791);
	dataBufferOut_long(4776) <= dataBufferIn_long( 792);
	dataBufferOut_long(5519) <= dataBufferIn_long( 793);
	dataBufferOut_long( 118) <= dataBufferIn_long( 794);
	dataBufferOut_long( 861) <= dataBufferIn_long( 795);
	dataBufferOut_long(1604) <= dataBufferIn_long( 796);
	dataBufferOut_long(2347) <= dataBufferIn_long( 797);
	dataBufferOut_long(3090) <= dataBufferIn_long( 798);
	dataBufferOut_long(3833) <= dataBufferIn_long( 799);
	dataBufferOut_long(4576) <= dataBufferIn_long( 800);
	dataBufferOut_long(5319) <= dataBufferIn_long( 801);
	dataBufferOut_long(6062) <= dataBufferIn_long( 802);
	dataBufferOut_long( 661) <= dataBufferIn_long( 803);
	dataBufferOut_long(1404) <= dataBufferIn_long( 804);
	dataBufferOut_long(2147) <= dataBufferIn_long( 805);
	dataBufferOut_long(2890) <= dataBufferIn_long( 806);
	dataBufferOut_long(3633) <= dataBufferIn_long( 807);
	dataBufferOut_long(4376) <= dataBufferIn_long( 808);
	dataBufferOut_long(5119) <= dataBufferIn_long( 809);
	dataBufferOut_long(5862) <= dataBufferIn_long( 810);
	dataBufferOut_long( 461) <= dataBufferIn_long( 811);
	dataBufferOut_long(1204) <= dataBufferIn_long( 812);
	dataBufferOut_long(1947) <= dataBufferIn_long( 813);
	dataBufferOut_long(2690) <= dataBufferIn_long( 814);
	dataBufferOut_long(3433) <= dataBufferIn_long( 815);
	dataBufferOut_long(4176) <= dataBufferIn_long( 816);
	dataBufferOut_long(4919) <= dataBufferIn_long( 817);
	dataBufferOut_long(5662) <= dataBufferIn_long( 818);
	dataBufferOut_long( 261) <= dataBufferIn_long( 819);
	dataBufferOut_long(1004) <= dataBufferIn_long( 820);
	dataBufferOut_long(1747) <= dataBufferIn_long( 821);
	dataBufferOut_long(2490) <= dataBufferIn_long( 822);
	dataBufferOut_long(3233) <= dataBufferIn_long( 823);
	dataBufferOut_long(3976) <= dataBufferIn_long( 824);
	dataBufferOut_long(4719) <= dataBufferIn_long( 825);
	dataBufferOut_long(5462) <= dataBufferIn_long( 826);
	dataBufferOut_long(  61) <= dataBufferIn_long( 827);
	dataBufferOut_long( 804) <= dataBufferIn_long( 828);
	dataBufferOut_long(1547) <= dataBufferIn_long( 829);
	dataBufferOut_long(2290) <= dataBufferIn_long( 830);
	dataBufferOut_long(3033) <= dataBufferIn_long( 831);
	dataBufferOut_long(3776) <= dataBufferIn_long( 832);
	dataBufferOut_long(4519) <= dataBufferIn_long( 833);
	dataBufferOut_long(5262) <= dataBufferIn_long( 834);
	dataBufferOut_long(6005) <= dataBufferIn_long( 835);
	dataBufferOut_long( 604) <= dataBufferIn_long( 836);
	dataBufferOut_long(1347) <= dataBufferIn_long( 837);
	dataBufferOut_long(2090) <= dataBufferIn_long( 838);
	dataBufferOut_long(2833) <= dataBufferIn_long( 839);
	dataBufferOut_long(3576) <= dataBufferIn_long( 840);
	dataBufferOut_long(4319) <= dataBufferIn_long( 841);
	dataBufferOut_long(5062) <= dataBufferIn_long( 842);
	dataBufferOut_long(5805) <= dataBufferIn_long( 843);
	dataBufferOut_long( 404) <= dataBufferIn_long( 844);
	dataBufferOut_long(1147) <= dataBufferIn_long( 845);
	dataBufferOut_long(1890) <= dataBufferIn_long( 846);
	dataBufferOut_long(2633) <= dataBufferIn_long( 847);
	dataBufferOut_long(3376) <= dataBufferIn_long( 848);
	dataBufferOut_long(4119) <= dataBufferIn_long( 849);
	dataBufferOut_long(4862) <= dataBufferIn_long( 850);
	dataBufferOut_long(5605) <= dataBufferIn_long( 851);
	dataBufferOut_long( 204) <= dataBufferIn_long( 852);
	dataBufferOut_long( 947) <= dataBufferIn_long( 853);
	dataBufferOut_long(1690) <= dataBufferIn_long( 854);
	dataBufferOut_long(2433) <= dataBufferIn_long( 855);
	dataBufferOut_long(3176) <= dataBufferIn_long( 856);
	dataBufferOut_long(3919) <= dataBufferIn_long( 857);
	dataBufferOut_long(4662) <= dataBufferIn_long( 858);
	dataBufferOut_long(5405) <= dataBufferIn_long( 859);
	dataBufferOut_long(   4) <= dataBufferIn_long( 860);
	dataBufferOut_long( 747) <= dataBufferIn_long( 861);
	dataBufferOut_long(1490) <= dataBufferIn_long( 862);
	dataBufferOut_long(2233) <= dataBufferIn_long( 863);
	dataBufferOut_long(2976) <= dataBufferIn_long( 864);
	dataBufferOut_long(3719) <= dataBufferIn_long( 865);
	dataBufferOut_long(4462) <= dataBufferIn_long( 866);
	dataBufferOut_long(5205) <= dataBufferIn_long( 867);
	dataBufferOut_long(5948) <= dataBufferIn_long( 868);
	dataBufferOut_long( 547) <= dataBufferIn_long( 869);
	dataBufferOut_long(1290) <= dataBufferIn_long( 870);
	dataBufferOut_long(2033) <= dataBufferIn_long( 871);
	dataBufferOut_long(2776) <= dataBufferIn_long( 872);
	dataBufferOut_long(3519) <= dataBufferIn_long( 873);
	dataBufferOut_long(4262) <= dataBufferIn_long( 874);
	dataBufferOut_long(5005) <= dataBufferIn_long( 875);
	dataBufferOut_long(5748) <= dataBufferIn_long( 876);
	dataBufferOut_long( 347) <= dataBufferIn_long( 877);
	dataBufferOut_long(1090) <= dataBufferIn_long( 878);
	dataBufferOut_long(1833) <= dataBufferIn_long( 879);
	dataBufferOut_long(2576) <= dataBufferIn_long( 880);
	dataBufferOut_long(3319) <= dataBufferIn_long( 881);
	dataBufferOut_long(4062) <= dataBufferIn_long( 882);
	dataBufferOut_long(4805) <= dataBufferIn_long( 883);
	dataBufferOut_long(5548) <= dataBufferIn_long( 884);
	dataBufferOut_long( 147) <= dataBufferIn_long( 885);
	dataBufferOut_long( 890) <= dataBufferIn_long( 886);
	dataBufferOut_long(1633) <= dataBufferIn_long( 887);
	dataBufferOut_long(2376) <= dataBufferIn_long( 888);
	dataBufferOut_long(3119) <= dataBufferIn_long( 889);
	dataBufferOut_long(3862) <= dataBufferIn_long( 890);
	dataBufferOut_long(4605) <= dataBufferIn_long( 891);
	dataBufferOut_long(5348) <= dataBufferIn_long( 892);
	dataBufferOut_long(6091) <= dataBufferIn_long( 893);
	dataBufferOut_long( 690) <= dataBufferIn_long( 894);
	dataBufferOut_long(1433) <= dataBufferIn_long( 895);
	dataBufferOut_long(2176) <= dataBufferIn_long( 896);
	dataBufferOut_long(2919) <= dataBufferIn_long( 897);
	dataBufferOut_long(3662) <= dataBufferIn_long( 898);
	dataBufferOut_long(4405) <= dataBufferIn_long( 899);
	dataBufferOut_long(5148) <= dataBufferIn_long( 900);
	dataBufferOut_long(5891) <= dataBufferIn_long( 901);
	dataBufferOut_long( 490) <= dataBufferIn_long( 902);
	dataBufferOut_long(1233) <= dataBufferIn_long( 903);
	dataBufferOut_long(1976) <= dataBufferIn_long( 904);
	dataBufferOut_long(2719) <= dataBufferIn_long( 905);
	dataBufferOut_long(3462) <= dataBufferIn_long( 906);
	dataBufferOut_long(4205) <= dataBufferIn_long( 907);
	dataBufferOut_long(4948) <= dataBufferIn_long( 908);
	dataBufferOut_long(5691) <= dataBufferIn_long( 909);
	dataBufferOut_long( 290) <= dataBufferIn_long( 910);
	dataBufferOut_long(1033) <= dataBufferIn_long( 911);
	dataBufferOut_long(1776) <= dataBufferIn_long( 912);
	dataBufferOut_long(2519) <= dataBufferIn_long( 913);
	dataBufferOut_long(3262) <= dataBufferIn_long( 914);
	dataBufferOut_long(4005) <= dataBufferIn_long( 915);
	dataBufferOut_long(4748) <= dataBufferIn_long( 916);
	dataBufferOut_long(5491) <= dataBufferIn_long( 917);
	dataBufferOut_long(  90) <= dataBufferIn_long( 918);
	dataBufferOut_long( 833) <= dataBufferIn_long( 919);
	dataBufferOut_long(1576) <= dataBufferIn_long( 920);
	dataBufferOut_long(2319) <= dataBufferIn_long( 921);
	dataBufferOut_long(3062) <= dataBufferIn_long( 922);
	dataBufferOut_long(3805) <= dataBufferIn_long( 923);
	dataBufferOut_long(4548) <= dataBufferIn_long( 924);
	dataBufferOut_long(5291) <= dataBufferIn_long( 925);
	dataBufferOut_long(6034) <= dataBufferIn_long( 926);
	dataBufferOut_long( 633) <= dataBufferIn_long( 927);
	dataBufferOut_long(1376) <= dataBufferIn_long( 928);
	dataBufferOut_long(2119) <= dataBufferIn_long( 929);
	dataBufferOut_long(2862) <= dataBufferIn_long( 930);
	dataBufferOut_long(3605) <= dataBufferIn_long( 931);
	dataBufferOut_long(4348) <= dataBufferIn_long( 932);
	dataBufferOut_long(5091) <= dataBufferIn_long( 933);
	dataBufferOut_long(5834) <= dataBufferIn_long( 934);
	dataBufferOut_long( 433) <= dataBufferIn_long( 935);
	dataBufferOut_long(1176) <= dataBufferIn_long( 936);
	dataBufferOut_long(1919) <= dataBufferIn_long( 937);
	dataBufferOut_long(2662) <= dataBufferIn_long( 938);
	dataBufferOut_long(3405) <= dataBufferIn_long( 939);
	dataBufferOut_long(4148) <= dataBufferIn_long( 940);
	dataBufferOut_long(4891) <= dataBufferIn_long( 941);
	dataBufferOut_long(5634) <= dataBufferIn_long( 942);
	dataBufferOut_long( 233) <= dataBufferIn_long( 943);
	dataBufferOut_long( 976) <= dataBufferIn_long( 944);
	dataBufferOut_long(1719) <= dataBufferIn_long( 945);
	dataBufferOut_long(2462) <= dataBufferIn_long( 946);
	dataBufferOut_long(3205) <= dataBufferIn_long( 947);
	dataBufferOut_long(3948) <= dataBufferIn_long( 948);
	dataBufferOut_long(4691) <= dataBufferIn_long( 949);
	dataBufferOut_long(5434) <= dataBufferIn_long( 950);
	dataBufferOut_long(  33) <= dataBufferIn_long( 951);
	dataBufferOut_long( 776) <= dataBufferIn_long( 952);
	dataBufferOut_long(1519) <= dataBufferIn_long( 953);
	dataBufferOut_long(2262) <= dataBufferIn_long( 954);
	dataBufferOut_long(3005) <= dataBufferIn_long( 955);
	dataBufferOut_long(3748) <= dataBufferIn_long( 956);
	dataBufferOut_long(4491) <= dataBufferIn_long( 957);
	dataBufferOut_long(5234) <= dataBufferIn_long( 958);
	dataBufferOut_long(5977) <= dataBufferIn_long( 959);
	dataBufferOut_long( 576) <= dataBufferIn_long( 960);
	dataBufferOut_long(1319) <= dataBufferIn_long( 961);
	dataBufferOut_long(2062) <= dataBufferIn_long( 962);
	dataBufferOut_long(2805) <= dataBufferIn_long( 963);
	dataBufferOut_long(3548) <= dataBufferIn_long( 964);
	dataBufferOut_long(4291) <= dataBufferIn_long( 965);
	dataBufferOut_long(5034) <= dataBufferIn_long( 966);
	dataBufferOut_long(5777) <= dataBufferIn_long( 967);
	dataBufferOut_long( 376) <= dataBufferIn_long( 968);
	dataBufferOut_long(1119) <= dataBufferIn_long( 969);
	dataBufferOut_long(1862) <= dataBufferIn_long( 970);
	dataBufferOut_long(2605) <= dataBufferIn_long( 971);
	dataBufferOut_long(3348) <= dataBufferIn_long( 972);
	dataBufferOut_long(4091) <= dataBufferIn_long( 973);
	dataBufferOut_long(4834) <= dataBufferIn_long( 974);
	dataBufferOut_long(5577) <= dataBufferIn_long( 975);
	dataBufferOut_long( 176) <= dataBufferIn_long( 976);
	dataBufferOut_long( 919) <= dataBufferIn_long( 977);
	dataBufferOut_long(1662) <= dataBufferIn_long( 978);
	dataBufferOut_long(2405) <= dataBufferIn_long( 979);
	dataBufferOut_long(3148) <= dataBufferIn_long( 980);
	dataBufferOut_long(3891) <= dataBufferIn_long( 981);
	dataBufferOut_long(4634) <= dataBufferIn_long( 982);
	dataBufferOut_long(5377) <= dataBufferIn_long( 983);
	dataBufferOut_long(6120) <= dataBufferIn_long( 984);
	dataBufferOut_long( 719) <= dataBufferIn_long( 985);
	dataBufferOut_long(1462) <= dataBufferIn_long( 986);
	dataBufferOut_long(2205) <= dataBufferIn_long( 987);
	dataBufferOut_long(2948) <= dataBufferIn_long( 988);
	dataBufferOut_long(3691) <= dataBufferIn_long( 989);
	dataBufferOut_long(4434) <= dataBufferIn_long( 990);
	dataBufferOut_long(5177) <= dataBufferIn_long( 991);
	dataBufferOut_long(5920) <= dataBufferIn_long( 992);
	dataBufferOut_long( 519) <= dataBufferIn_long( 993);
	dataBufferOut_long(1262) <= dataBufferIn_long( 994);
	dataBufferOut_long(2005) <= dataBufferIn_long( 995);
	dataBufferOut_long(2748) <= dataBufferIn_long( 996);
	dataBufferOut_long(3491) <= dataBufferIn_long( 997);
	dataBufferOut_long(4234) <= dataBufferIn_long( 998);
	dataBufferOut_long(4977) <= dataBufferIn_long( 999);
	dataBufferOut_long(5720) <= dataBufferIn_long(1000);
	dataBufferOut_long( 319) <= dataBufferIn_long(1001);
	dataBufferOut_long(1062) <= dataBufferIn_long(1002);
	dataBufferOut_long(1805) <= dataBufferIn_long(1003);
	dataBufferOut_long(2548) <= dataBufferIn_long(1004);
	dataBufferOut_long(3291) <= dataBufferIn_long(1005);
	dataBufferOut_long(4034) <= dataBufferIn_long(1006);
	dataBufferOut_long(4777) <= dataBufferIn_long(1007);
	dataBufferOut_long(5520) <= dataBufferIn_long(1008);
	dataBufferOut_long( 119) <= dataBufferIn_long(1009);
	dataBufferOut_long( 862) <= dataBufferIn_long(1010);
	dataBufferOut_long(1605) <= dataBufferIn_long(1011);
	dataBufferOut_long(2348) <= dataBufferIn_long(1012);
	dataBufferOut_long(3091) <= dataBufferIn_long(1013);
	dataBufferOut_long(3834) <= dataBufferIn_long(1014);
	dataBufferOut_long(4577) <= dataBufferIn_long(1015);
	dataBufferOut_long(5320) <= dataBufferIn_long(1016);
	dataBufferOut_long(6063) <= dataBufferIn_long(1017);
	dataBufferOut_long( 662) <= dataBufferIn_long(1018);
	dataBufferOut_long(1405) <= dataBufferIn_long(1019);
	dataBufferOut_long(2148) <= dataBufferIn_long(1020);
	dataBufferOut_long(2891) <= dataBufferIn_long(1021);
	dataBufferOut_long(3634) <= dataBufferIn_long(1022);
	dataBufferOut_long(4377) <= dataBufferIn_long(1023);
	dataBufferOut_long(5120) <= dataBufferIn_long(1024);
	dataBufferOut_long(5863) <= dataBufferIn_long(1025);
	dataBufferOut_long( 462) <= dataBufferIn_long(1026);
	dataBufferOut_long(1205) <= dataBufferIn_long(1027);
	dataBufferOut_long(1948) <= dataBufferIn_long(1028);
	dataBufferOut_long(2691) <= dataBufferIn_long(1029);
	dataBufferOut_long(3434) <= dataBufferIn_long(1030);
	dataBufferOut_long(4177) <= dataBufferIn_long(1031);
	dataBufferOut_long(4920) <= dataBufferIn_long(1032);
	dataBufferOut_long(5663) <= dataBufferIn_long(1033);
	dataBufferOut_long( 262) <= dataBufferIn_long(1034);
	dataBufferOut_long(1005) <= dataBufferIn_long(1035);
	dataBufferOut_long(1748) <= dataBufferIn_long(1036);
	dataBufferOut_long(2491) <= dataBufferIn_long(1037);
	dataBufferOut_long(3234) <= dataBufferIn_long(1038);
	dataBufferOut_long(3977) <= dataBufferIn_long(1039);
	dataBufferOut_long(4720) <= dataBufferIn_long(1040);
	dataBufferOut_long(5463) <= dataBufferIn_long(1041);
	dataBufferOut_long(  62) <= dataBufferIn_long(1042);
	dataBufferOut_long( 805) <= dataBufferIn_long(1043);
	dataBufferOut_long(1548) <= dataBufferIn_long(1044);
	dataBufferOut_long(2291) <= dataBufferIn_long(1045);
	dataBufferOut_long(3034) <= dataBufferIn_long(1046);
	dataBufferOut_long(3777) <= dataBufferIn_long(1047);
	dataBufferOut_long(4520) <= dataBufferIn_long(1048);
	dataBufferOut_long(5263) <= dataBufferIn_long(1049);
	dataBufferOut_long(6006) <= dataBufferIn_long(1050);
	dataBufferOut_long( 605) <= dataBufferIn_long(1051);
	dataBufferOut_long(1348) <= dataBufferIn_long(1052);
	dataBufferOut_long(2091) <= dataBufferIn_long(1053);
	dataBufferOut_long(2834) <= dataBufferIn_long(1054);
	dataBufferOut_long(3577) <= dataBufferIn_long(1055);
	dataBufferOut_long(4320) <= dataBufferIn_long(1056);
	dataBufferOut_long(5063) <= dataBufferIn_long(1057);
	dataBufferOut_long(5806) <= dataBufferIn_long(1058);
	dataBufferOut_long( 405) <= dataBufferIn_long(1059);
	dataBufferOut_long(1148) <= dataBufferIn_long(1060);
	dataBufferOut_long(1891) <= dataBufferIn_long(1061);
	dataBufferOut_long(2634) <= dataBufferIn_long(1062);
	dataBufferOut_long(3377) <= dataBufferIn_long(1063);
	dataBufferOut_long(4120) <= dataBufferIn_long(1064);
	dataBufferOut_long(4863) <= dataBufferIn_long(1065);
	dataBufferOut_long(5606) <= dataBufferIn_long(1066);
	dataBufferOut_long( 205) <= dataBufferIn_long(1067);
	dataBufferOut_long( 948) <= dataBufferIn_long(1068);
	dataBufferOut_long(1691) <= dataBufferIn_long(1069);
	dataBufferOut_long(2434) <= dataBufferIn_long(1070);
	dataBufferOut_long(3177) <= dataBufferIn_long(1071);
	dataBufferOut_long(3920) <= dataBufferIn_long(1072);
	dataBufferOut_long(4663) <= dataBufferIn_long(1073);
	dataBufferOut_long(5406) <= dataBufferIn_long(1074);
	dataBufferOut_long(   5) <= dataBufferIn_long(1075);
	dataBufferOut_long( 748) <= dataBufferIn_long(1076);
	dataBufferOut_long(1491) <= dataBufferIn_long(1077);
	dataBufferOut_long(2234) <= dataBufferIn_long(1078);
	dataBufferOut_long(2977) <= dataBufferIn_long(1079);
	dataBufferOut_long(3720) <= dataBufferIn_long(1080);
	dataBufferOut_long(4463) <= dataBufferIn_long(1081);
	dataBufferOut_long(5206) <= dataBufferIn_long(1082);
	dataBufferOut_long(5949) <= dataBufferIn_long(1083);
	dataBufferOut_long( 548) <= dataBufferIn_long(1084);
	dataBufferOut_long(1291) <= dataBufferIn_long(1085);
	dataBufferOut_long(2034) <= dataBufferIn_long(1086);
	dataBufferOut_long(2777) <= dataBufferIn_long(1087);
	dataBufferOut_long(3520) <= dataBufferIn_long(1088);
	dataBufferOut_long(4263) <= dataBufferIn_long(1089);
	dataBufferOut_long(5006) <= dataBufferIn_long(1090);
	dataBufferOut_long(5749) <= dataBufferIn_long(1091);
	dataBufferOut_long( 348) <= dataBufferIn_long(1092);
	dataBufferOut_long(1091) <= dataBufferIn_long(1093);
	dataBufferOut_long(1834) <= dataBufferIn_long(1094);
	dataBufferOut_long(2577) <= dataBufferIn_long(1095);
	dataBufferOut_long(3320) <= dataBufferIn_long(1096);
	dataBufferOut_long(4063) <= dataBufferIn_long(1097);
	dataBufferOut_long(4806) <= dataBufferIn_long(1098);
	dataBufferOut_long(5549) <= dataBufferIn_long(1099);
	dataBufferOut_long( 148) <= dataBufferIn_long(1100);
	dataBufferOut_long( 891) <= dataBufferIn_long(1101);
	dataBufferOut_long(1634) <= dataBufferIn_long(1102);
	dataBufferOut_long(2377) <= dataBufferIn_long(1103);
	dataBufferOut_long(3120) <= dataBufferIn_long(1104);
	dataBufferOut_long(3863) <= dataBufferIn_long(1105);
	dataBufferOut_long(4606) <= dataBufferIn_long(1106);
	dataBufferOut_long(5349) <= dataBufferIn_long(1107);
	dataBufferOut_long(6092) <= dataBufferIn_long(1108);
	dataBufferOut_long( 691) <= dataBufferIn_long(1109);
	dataBufferOut_long(1434) <= dataBufferIn_long(1110);
	dataBufferOut_long(2177) <= dataBufferIn_long(1111);
	dataBufferOut_long(2920) <= dataBufferIn_long(1112);
	dataBufferOut_long(3663) <= dataBufferIn_long(1113);
	dataBufferOut_long(4406) <= dataBufferIn_long(1114);
	dataBufferOut_long(5149) <= dataBufferIn_long(1115);
	dataBufferOut_long(5892) <= dataBufferIn_long(1116);
	dataBufferOut_long( 491) <= dataBufferIn_long(1117);
	dataBufferOut_long(1234) <= dataBufferIn_long(1118);
	dataBufferOut_long(1977) <= dataBufferIn_long(1119);
	dataBufferOut_long(2720) <= dataBufferIn_long(1120);
	dataBufferOut_long(3463) <= dataBufferIn_long(1121);
	dataBufferOut_long(4206) <= dataBufferIn_long(1122);
	dataBufferOut_long(4949) <= dataBufferIn_long(1123);
	dataBufferOut_long(5692) <= dataBufferIn_long(1124);
	dataBufferOut_long( 291) <= dataBufferIn_long(1125);
	dataBufferOut_long(1034) <= dataBufferIn_long(1126);
	dataBufferOut_long(1777) <= dataBufferIn_long(1127);
	dataBufferOut_long(2520) <= dataBufferIn_long(1128);
	dataBufferOut_long(3263) <= dataBufferIn_long(1129);
	dataBufferOut_long(4006) <= dataBufferIn_long(1130);
	dataBufferOut_long(4749) <= dataBufferIn_long(1131);
	dataBufferOut_long(5492) <= dataBufferIn_long(1132);
	dataBufferOut_long(  91) <= dataBufferIn_long(1133);
	dataBufferOut_long( 834) <= dataBufferIn_long(1134);
	dataBufferOut_long(1577) <= dataBufferIn_long(1135);
	dataBufferOut_long(2320) <= dataBufferIn_long(1136);
	dataBufferOut_long(3063) <= dataBufferIn_long(1137);
	dataBufferOut_long(3806) <= dataBufferIn_long(1138);
	dataBufferOut_long(4549) <= dataBufferIn_long(1139);
	dataBufferOut_long(5292) <= dataBufferIn_long(1140);
	dataBufferOut_long(6035) <= dataBufferIn_long(1141);
	dataBufferOut_long( 634) <= dataBufferIn_long(1142);
	dataBufferOut_long(1377) <= dataBufferIn_long(1143);
	dataBufferOut_long(2120) <= dataBufferIn_long(1144);
	dataBufferOut_long(2863) <= dataBufferIn_long(1145);
	dataBufferOut_long(3606) <= dataBufferIn_long(1146);
	dataBufferOut_long(4349) <= dataBufferIn_long(1147);
	dataBufferOut_long(5092) <= dataBufferIn_long(1148);
	dataBufferOut_long(5835) <= dataBufferIn_long(1149);
	dataBufferOut_long( 434) <= dataBufferIn_long(1150);
	dataBufferOut_long(1177) <= dataBufferIn_long(1151);
	dataBufferOut_long(1920) <= dataBufferIn_long(1152);
	dataBufferOut_long(2663) <= dataBufferIn_long(1153);
	dataBufferOut_long(3406) <= dataBufferIn_long(1154);
	dataBufferOut_long(4149) <= dataBufferIn_long(1155);
	dataBufferOut_long(4892) <= dataBufferIn_long(1156);
	dataBufferOut_long(5635) <= dataBufferIn_long(1157);
	dataBufferOut_long( 234) <= dataBufferIn_long(1158);
	dataBufferOut_long( 977) <= dataBufferIn_long(1159);
	dataBufferOut_long(1720) <= dataBufferIn_long(1160);
	dataBufferOut_long(2463) <= dataBufferIn_long(1161);
	dataBufferOut_long(3206) <= dataBufferIn_long(1162);
	dataBufferOut_long(3949) <= dataBufferIn_long(1163);
	dataBufferOut_long(4692) <= dataBufferIn_long(1164);
	dataBufferOut_long(5435) <= dataBufferIn_long(1165);
	dataBufferOut_long(  34) <= dataBufferIn_long(1166);
	dataBufferOut_long( 777) <= dataBufferIn_long(1167);
	dataBufferOut_long(1520) <= dataBufferIn_long(1168);
	dataBufferOut_long(2263) <= dataBufferIn_long(1169);
	dataBufferOut_long(3006) <= dataBufferIn_long(1170);
	dataBufferOut_long(3749) <= dataBufferIn_long(1171);
	dataBufferOut_long(4492) <= dataBufferIn_long(1172);
	dataBufferOut_long(5235) <= dataBufferIn_long(1173);
	dataBufferOut_long(5978) <= dataBufferIn_long(1174);
	dataBufferOut_long( 577) <= dataBufferIn_long(1175);
	dataBufferOut_long(1320) <= dataBufferIn_long(1176);
	dataBufferOut_long(2063) <= dataBufferIn_long(1177);
	dataBufferOut_long(2806) <= dataBufferIn_long(1178);
	dataBufferOut_long(3549) <= dataBufferIn_long(1179);
	dataBufferOut_long(4292) <= dataBufferIn_long(1180);
	dataBufferOut_long(5035) <= dataBufferIn_long(1181);
	dataBufferOut_long(5778) <= dataBufferIn_long(1182);
	dataBufferOut_long( 377) <= dataBufferIn_long(1183);
	dataBufferOut_long(1120) <= dataBufferIn_long(1184);
	dataBufferOut_long(1863) <= dataBufferIn_long(1185);
	dataBufferOut_long(2606) <= dataBufferIn_long(1186);
	dataBufferOut_long(3349) <= dataBufferIn_long(1187);
	dataBufferOut_long(4092) <= dataBufferIn_long(1188);
	dataBufferOut_long(4835) <= dataBufferIn_long(1189);
	dataBufferOut_long(5578) <= dataBufferIn_long(1190);
	dataBufferOut_long( 177) <= dataBufferIn_long(1191);
	dataBufferOut_long( 920) <= dataBufferIn_long(1192);
	dataBufferOut_long(1663) <= dataBufferIn_long(1193);
	dataBufferOut_long(2406) <= dataBufferIn_long(1194);
	dataBufferOut_long(3149) <= dataBufferIn_long(1195);
	dataBufferOut_long(3892) <= dataBufferIn_long(1196);
	dataBufferOut_long(4635) <= dataBufferIn_long(1197);
	dataBufferOut_long(5378) <= dataBufferIn_long(1198);
	dataBufferOut_long(6121) <= dataBufferIn_long(1199);
	dataBufferOut_long( 720) <= dataBufferIn_long(1200);
	dataBufferOut_long(1463) <= dataBufferIn_long(1201);
	dataBufferOut_long(2206) <= dataBufferIn_long(1202);
	dataBufferOut_long(2949) <= dataBufferIn_long(1203);
	dataBufferOut_long(3692) <= dataBufferIn_long(1204);
	dataBufferOut_long(4435) <= dataBufferIn_long(1205);
	dataBufferOut_long(5178) <= dataBufferIn_long(1206);
	dataBufferOut_long(5921) <= dataBufferIn_long(1207);
	dataBufferOut_long( 520) <= dataBufferIn_long(1208);
	dataBufferOut_long(1263) <= dataBufferIn_long(1209);
	dataBufferOut_long(2006) <= dataBufferIn_long(1210);
	dataBufferOut_long(2749) <= dataBufferIn_long(1211);
	dataBufferOut_long(3492) <= dataBufferIn_long(1212);
	dataBufferOut_long(4235) <= dataBufferIn_long(1213);
	dataBufferOut_long(4978) <= dataBufferIn_long(1214);
	dataBufferOut_long(5721) <= dataBufferIn_long(1215);
	dataBufferOut_long( 320) <= dataBufferIn_long(1216);
	dataBufferOut_long(1063) <= dataBufferIn_long(1217);
	dataBufferOut_long(1806) <= dataBufferIn_long(1218);
	dataBufferOut_long(2549) <= dataBufferIn_long(1219);
	dataBufferOut_long(3292) <= dataBufferIn_long(1220);
	dataBufferOut_long(4035) <= dataBufferIn_long(1221);
	dataBufferOut_long(4778) <= dataBufferIn_long(1222);
	dataBufferOut_long(5521) <= dataBufferIn_long(1223);
	dataBufferOut_long( 120) <= dataBufferIn_long(1224);
	dataBufferOut_long( 863) <= dataBufferIn_long(1225);
	dataBufferOut_long(1606) <= dataBufferIn_long(1226);
	dataBufferOut_long(2349) <= dataBufferIn_long(1227);
	dataBufferOut_long(3092) <= dataBufferIn_long(1228);
	dataBufferOut_long(3835) <= dataBufferIn_long(1229);
	dataBufferOut_long(4578) <= dataBufferIn_long(1230);
	dataBufferOut_long(5321) <= dataBufferIn_long(1231);
	dataBufferOut_long(6064) <= dataBufferIn_long(1232);
	dataBufferOut_long( 663) <= dataBufferIn_long(1233);
	dataBufferOut_long(1406) <= dataBufferIn_long(1234);
	dataBufferOut_long(2149) <= dataBufferIn_long(1235);
	dataBufferOut_long(2892) <= dataBufferIn_long(1236);
	dataBufferOut_long(3635) <= dataBufferIn_long(1237);
	dataBufferOut_long(4378) <= dataBufferIn_long(1238);
	dataBufferOut_long(5121) <= dataBufferIn_long(1239);
	dataBufferOut_long(5864) <= dataBufferIn_long(1240);
	dataBufferOut_long( 463) <= dataBufferIn_long(1241);
	dataBufferOut_long(1206) <= dataBufferIn_long(1242);
	dataBufferOut_long(1949) <= dataBufferIn_long(1243);
	dataBufferOut_long(2692) <= dataBufferIn_long(1244);
	dataBufferOut_long(3435) <= dataBufferIn_long(1245);
	dataBufferOut_long(4178) <= dataBufferIn_long(1246);
	dataBufferOut_long(4921) <= dataBufferIn_long(1247);
	dataBufferOut_long(5664) <= dataBufferIn_long(1248);
	dataBufferOut_long( 263) <= dataBufferIn_long(1249);
	dataBufferOut_long(1006) <= dataBufferIn_long(1250);
	dataBufferOut_long(1749) <= dataBufferIn_long(1251);
	dataBufferOut_long(2492) <= dataBufferIn_long(1252);
	dataBufferOut_long(3235) <= dataBufferIn_long(1253);
	dataBufferOut_long(3978) <= dataBufferIn_long(1254);
	dataBufferOut_long(4721) <= dataBufferIn_long(1255);
	dataBufferOut_long(5464) <= dataBufferIn_long(1256);
	dataBufferOut_long(  63) <= dataBufferIn_long(1257);
	dataBufferOut_long( 806) <= dataBufferIn_long(1258);
	dataBufferOut_long(1549) <= dataBufferIn_long(1259);
	dataBufferOut_long(2292) <= dataBufferIn_long(1260);
	dataBufferOut_long(3035) <= dataBufferIn_long(1261);
	dataBufferOut_long(3778) <= dataBufferIn_long(1262);
	dataBufferOut_long(4521) <= dataBufferIn_long(1263);
	dataBufferOut_long(5264) <= dataBufferIn_long(1264);
	dataBufferOut_long(6007) <= dataBufferIn_long(1265);
	dataBufferOut_long( 606) <= dataBufferIn_long(1266);
	dataBufferOut_long(1349) <= dataBufferIn_long(1267);
	dataBufferOut_long(2092) <= dataBufferIn_long(1268);
	dataBufferOut_long(2835) <= dataBufferIn_long(1269);
	dataBufferOut_long(3578) <= dataBufferIn_long(1270);
	dataBufferOut_long(4321) <= dataBufferIn_long(1271);
	dataBufferOut_long(5064) <= dataBufferIn_long(1272);
	dataBufferOut_long(5807) <= dataBufferIn_long(1273);
	dataBufferOut_long( 406) <= dataBufferIn_long(1274);
	dataBufferOut_long(1149) <= dataBufferIn_long(1275);
	dataBufferOut_long(1892) <= dataBufferIn_long(1276);
	dataBufferOut_long(2635) <= dataBufferIn_long(1277);
	dataBufferOut_long(3378) <= dataBufferIn_long(1278);
	dataBufferOut_long(4121) <= dataBufferIn_long(1279);
	dataBufferOut_long(4864) <= dataBufferIn_long(1280);
	dataBufferOut_long(5607) <= dataBufferIn_long(1281);
	dataBufferOut_long( 206) <= dataBufferIn_long(1282);
	dataBufferOut_long( 949) <= dataBufferIn_long(1283);
	dataBufferOut_long(1692) <= dataBufferIn_long(1284);
	dataBufferOut_long(2435) <= dataBufferIn_long(1285);
	dataBufferOut_long(3178) <= dataBufferIn_long(1286);
	dataBufferOut_long(3921) <= dataBufferIn_long(1287);
	dataBufferOut_long(4664) <= dataBufferIn_long(1288);
	dataBufferOut_long(5407) <= dataBufferIn_long(1289);
	dataBufferOut_long(   6) <= dataBufferIn_long(1290);
	dataBufferOut_long( 749) <= dataBufferIn_long(1291);
	dataBufferOut_long(1492) <= dataBufferIn_long(1292);
	dataBufferOut_long(2235) <= dataBufferIn_long(1293);
	dataBufferOut_long(2978) <= dataBufferIn_long(1294);
	dataBufferOut_long(3721) <= dataBufferIn_long(1295);
	dataBufferOut_long(4464) <= dataBufferIn_long(1296);
	dataBufferOut_long(5207) <= dataBufferIn_long(1297);
	dataBufferOut_long(5950) <= dataBufferIn_long(1298);
	dataBufferOut_long( 549) <= dataBufferIn_long(1299);
	dataBufferOut_long(1292) <= dataBufferIn_long(1300);
	dataBufferOut_long(2035) <= dataBufferIn_long(1301);
	dataBufferOut_long(2778) <= dataBufferIn_long(1302);
	dataBufferOut_long(3521) <= dataBufferIn_long(1303);
	dataBufferOut_long(4264) <= dataBufferIn_long(1304);
	dataBufferOut_long(5007) <= dataBufferIn_long(1305);
	dataBufferOut_long(5750) <= dataBufferIn_long(1306);
	dataBufferOut_long( 349) <= dataBufferIn_long(1307);
	dataBufferOut_long(1092) <= dataBufferIn_long(1308);
	dataBufferOut_long(1835) <= dataBufferIn_long(1309);
	dataBufferOut_long(2578) <= dataBufferIn_long(1310);
	dataBufferOut_long(3321) <= dataBufferIn_long(1311);
	dataBufferOut_long(4064) <= dataBufferIn_long(1312);
	dataBufferOut_long(4807) <= dataBufferIn_long(1313);
	dataBufferOut_long(5550) <= dataBufferIn_long(1314);
	dataBufferOut_long( 149) <= dataBufferIn_long(1315);
	dataBufferOut_long( 892) <= dataBufferIn_long(1316);
	dataBufferOut_long(1635) <= dataBufferIn_long(1317);
	dataBufferOut_long(2378) <= dataBufferIn_long(1318);
	dataBufferOut_long(3121) <= dataBufferIn_long(1319);
	dataBufferOut_long(3864) <= dataBufferIn_long(1320);
	dataBufferOut_long(4607) <= dataBufferIn_long(1321);
	dataBufferOut_long(5350) <= dataBufferIn_long(1322);
	dataBufferOut_long(6093) <= dataBufferIn_long(1323);
	dataBufferOut_long( 692) <= dataBufferIn_long(1324);
	dataBufferOut_long(1435) <= dataBufferIn_long(1325);
	dataBufferOut_long(2178) <= dataBufferIn_long(1326);
	dataBufferOut_long(2921) <= dataBufferIn_long(1327);
	dataBufferOut_long(3664) <= dataBufferIn_long(1328);
	dataBufferOut_long(4407) <= dataBufferIn_long(1329);
	dataBufferOut_long(5150) <= dataBufferIn_long(1330);
	dataBufferOut_long(5893) <= dataBufferIn_long(1331);
	dataBufferOut_long( 492) <= dataBufferIn_long(1332);
	dataBufferOut_long(1235) <= dataBufferIn_long(1333);
	dataBufferOut_long(1978) <= dataBufferIn_long(1334);
	dataBufferOut_long(2721) <= dataBufferIn_long(1335);
	dataBufferOut_long(3464) <= dataBufferIn_long(1336);
	dataBufferOut_long(4207) <= dataBufferIn_long(1337);
	dataBufferOut_long(4950) <= dataBufferIn_long(1338);
	dataBufferOut_long(5693) <= dataBufferIn_long(1339);
	dataBufferOut_long( 292) <= dataBufferIn_long(1340);
	dataBufferOut_long(1035) <= dataBufferIn_long(1341);
	dataBufferOut_long(1778) <= dataBufferIn_long(1342);
	dataBufferOut_long(2521) <= dataBufferIn_long(1343);
	dataBufferOut_long(3264) <= dataBufferIn_long(1344);
	dataBufferOut_long(4007) <= dataBufferIn_long(1345);
	dataBufferOut_long(4750) <= dataBufferIn_long(1346);
	dataBufferOut_long(5493) <= dataBufferIn_long(1347);
	dataBufferOut_long(  92) <= dataBufferIn_long(1348);
	dataBufferOut_long( 835) <= dataBufferIn_long(1349);
	dataBufferOut_long(1578) <= dataBufferIn_long(1350);
	dataBufferOut_long(2321) <= dataBufferIn_long(1351);
	dataBufferOut_long(3064) <= dataBufferIn_long(1352);
	dataBufferOut_long(3807) <= dataBufferIn_long(1353);
	dataBufferOut_long(4550) <= dataBufferIn_long(1354);
	dataBufferOut_long(5293) <= dataBufferIn_long(1355);
	dataBufferOut_long(6036) <= dataBufferIn_long(1356);
	dataBufferOut_long( 635) <= dataBufferIn_long(1357);
	dataBufferOut_long(1378) <= dataBufferIn_long(1358);
	dataBufferOut_long(2121) <= dataBufferIn_long(1359);
	dataBufferOut_long(2864) <= dataBufferIn_long(1360);
	dataBufferOut_long(3607) <= dataBufferIn_long(1361);
	dataBufferOut_long(4350) <= dataBufferIn_long(1362);
	dataBufferOut_long(5093) <= dataBufferIn_long(1363);
	dataBufferOut_long(5836) <= dataBufferIn_long(1364);
	dataBufferOut_long( 435) <= dataBufferIn_long(1365);
	dataBufferOut_long(1178) <= dataBufferIn_long(1366);
	dataBufferOut_long(1921) <= dataBufferIn_long(1367);
	dataBufferOut_long(2664) <= dataBufferIn_long(1368);
	dataBufferOut_long(3407) <= dataBufferIn_long(1369);
	dataBufferOut_long(4150) <= dataBufferIn_long(1370);
	dataBufferOut_long(4893) <= dataBufferIn_long(1371);
	dataBufferOut_long(5636) <= dataBufferIn_long(1372);
	dataBufferOut_long( 235) <= dataBufferIn_long(1373);
	dataBufferOut_long( 978) <= dataBufferIn_long(1374);
	dataBufferOut_long(1721) <= dataBufferIn_long(1375);
	dataBufferOut_long(2464) <= dataBufferIn_long(1376);
	dataBufferOut_long(3207) <= dataBufferIn_long(1377);
	dataBufferOut_long(3950) <= dataBufferIn_long(1378);
	dataBufferOut_long(4693) <= dataBufferIn_long(1379);
	dataBufferOut_long(5436) <= dataBufferIn_long(1380);
	dataBufferOut_long(  35) <= dataBufferIn_long(1381);
	dataBufferOut_long( 778) <= dataBufferIn_long(1382);
	dataBufferOut_long(1521) <= dataBufferIn_long(1383);
	dataBufferOut_long(2264) <= dataBufferIn_long(1384);
	dataBufferOut_long(3007) <= dataBufferIn_long(1385);
	dataBufferOut_long(3750) <= dataBufferIn_long(1386);
	dataBufferOut_long(4493) <= dataBufferIn_long(1387);
	dataBufferOut_long(5236) <= dataBufferIn_long(1388);
	dataBufferOut_long(5979) <= dataBufferIn_long(1389);
	dataBufferOut_long( 578) <= dataBufferIn_long(1390);
	dataBufferOut_long(1321) <= dataBufferIn_long(1391);
	dataBufferOut_long(2064) <= dataBufferIn_long(1392);
	dataBufferOut_long(2807) <= dataBufferIn_long(1393);
	dataBufferOut_long(3550) <= dataBufferIn_long(1394);
	dataBufferOut_long(4293) <= dataBufferIn_long(1395);
	dataBufferOut_long(5036) <= dataBufferIn_long(1396);
	dataBufferOut_long(5779) <= dataBufferIn_long(1397);
	dataBufferOut_long( 378) <= dataBufferIn_long(1398);
	dataBufferOut_long(1121) <= dataBufferIn_long(1399);
	dataBufferOut_long(1864) <= dataBufferIn_long(1400);
	dataBufferOut_long(2607) <= dataBufferIn_long(1401);
	dataBufferOut_long(3350) <= dataBufferIn_long(1402);
	dataBufferOut_long(4093) <= dataBufferIn_long(1403);
	dataBufferOut_long(4836) <= dataBufferIn_long(1404);
	dataBufferOut_long(5579) <= dataBufferIn_long(1405);
	dataBufferOut_long( 178) <= dataBufferIn_long(1406);
	dataBufferOut_long( 921) <= dataBufferIn_long(1407);
	dataBufferOut_long(1664) <= dataBufferIn_long(1408);
	dataBufferOut_long(2407) <= dataBufferIn_long(1409);
	dataBufferOut_long(3150) <= dataBufferIn_long(1410);
	dataBufferOut_long(3893) <= dataBufferIn_long(1411);
	dataBufferOut_long(4636) <= dataBufferIn_long(1412);
	dataBufferOut_long(5379) <= dataBufferIn_long(1413);
	dataBufferOut_long(6122) <= dataBufferIn_long(1414);
	dataBufferOut_long( 721) <= dataBufferIn_long(1415);
	dataBufferOut_long(1464) <= dataBufferIn_long(1416);
	dataBufferOut_long(2207) <= dataBufferIn_long(1417);
	dataBufferOut_long(2950) <= dataBufferIn_long(1418);
	dataBufferOut_long(3693) <= dataBufferIn_long(1419);
	dataBufferOut_long(4436) <= dataBufferIn_long(1420);
	dataBufferOut_long(5179) <= dataBufferIn_long(1421);
	dataBufferOut_long(5922) <= dataBufferIn_long(1422);
	dataBufferOut_long( 521) <= dataBufferIn_long(1423);
	dataBufferOut_long(1264) <= dataBufferIn_long(1424);
	dataBufferOut_long(2007) <= dataBufferIn_long(1425);
	dataBufferOut_long(2750) <= dataBufferIn_long(1426);
	dataBufferOut_long(3493) <= dataBufferIn_long(1427);
	dataBufferOut_long(4236) <= dataBufferIn_long(1428);
	dataBufferOut_long(4979) <= dataBufferIn_long(1429);
	dataBufferOut_long(5722) <= dataBufferIn_long(1430);
	dataBufferOut_long( 321) <= dataBufferIn_long(1431);
	dataBufferOut_long(1064) <= dataBufferIn_long(1432);
	dataBufferOut_long(1807) <= dataBufferIn_long(1433);
	dataBufferOut_long(2550) <= dataBufferIn_long(1434);
	dataBufferOut_long(3293) <= dataBufferIn_long(1435);
	dataBufferOut_long(4036) <= dataBufferIn_long(1436);
	dataBufferOut_long(4779) <= dataBufferIn_long(1437);
	dataBufferOut_long(5522) <= dataBufferIn_long(1438);
	dataBufferOut_long( 121) <= dataBufferIn_long(1439);
	dataBufferOut_long( 864) <= dataBufferIn_long(1440);
	dataBufferOut_long(1607) <= dataBufferIn_long(1441);
	dataBufferOut_long(2350) <= dataBufferIn_long(1442);
	dataBufferOut_long(3093) <= dataBufferIn_long(1443);
	dataBufferOut_long(3836) <= dataBufferIn_long(1444);
	dataBufferOut_long(4579) <= dataBufferIn_long(1445);
	dataBufferOut_long(5322) <= dataBufferIn_long(1446);
	dataBufferOut_long(6065) <= dataBufferIn_long(1447);
	dataBufferOut_long( 664) <= dataBufferIn_long(1448);
	dataBufferOut_long(1407) <= dataBufferIn_long(1449);
	dataBufferOut_long(2150) <= dataBufferIn_long(1450);
	dataBufferOut_long(2893) <= dataBufferIn_long(1451);
	dataBufferOut_long(3636) <= dataBufferIn_long(1452);
	dataBufferOut_long(4379) <= dataBufferIn_long(1453);
	dataBufferOut_long(5122) <= dataBufferIn_long(1454);
	dataBufferOut_long(5865) <= dataBufferIn_long(1455);
	dataBufferOut_long( 464) <= dataBufferIn_long(1456);
	dataBufferOut_long(1207) <= dataBufferIn_long(1457);
	dataBufferOut_long(1950) <= dataBufferIn_long(1458);
	dataBufferOut_long(2693) <= dataBufferIn_long(1459);
	dataBufferOut_long(3436) <= dataBufferIn_long(1460);
	dataBufferOut_long(4179) <= dataBufferIn_long(1461);
	dataBufferOut_long(4922) <= dataBufferIn_long(1462);
	dataBufferOut_long(5665) <= dataBufferIn_long(1463);
	dataBufferOut_long( 264) <= dataBufferIn_long(1464);
	dataBufferOut_long(1007) <= dataBufferIn_long(1465);
	dataBufferOut_long(1750) <= dataBufferIn_long(1466);
	dataBufferOut_long(2493) <= dataBufferIn_long(1467);
	dataBufferOut_long(3236) <= dataBufferIn_long(1468);
	dataBufferOut_long(3979) <= dataBufferIn_long(1469);
	dataBufferOut_long(4722) <= dataBufferIn_long(1470);
	dataBufferOut_long(5465) <= dataBufferIn_long(1471);
	dataBufferOut_long(  64) <= dataBufferIn_long(1472);
	dataBufferOut_long( 807) <= dataBufferIn_long(1473);
	dataBufferOut_long(1550) <= dataBufferIn_long(1474);
	dataBufferOut_long(2293) <= dataBufferIn_long(1475);
	dataBufferOut_long(3036) <= dataBufferIn_long(1476);
	dataBufferOut_long(3779) <= dataBufferIn_long(1477);
	dataBufferOut_long(4522) <= dataBufferIn_long(1478);
	dataBufferOut_long(5265) <= dataBufferIn_long(1479);
	dataBufferOut_long(6008) <= dataBufferIn_long(1480);
	dataBufferOut_long( 607) <= dataBufferIn_long(1481);
	dataBufferOut_long(1350) <= dataBufferIn_long(1482);
	dataBufferOut_long(2093) <= dataBufferIn_long(1483);
	dataBufferOut_long(2836) <= dataBufferIn_long(1484);
	dataBufferOut_long(3579) <= dataBufferIn_long(1485);
	dataBufferOut_long(4322) <= dataBufferIn_long(1486);
	dataBufferOut_long(5065) <= dataBufferIn_long(1487);
	dataBufferOut_long(5808) <= dataBufferIn_long(1488);
	dataBufferOut_long( 407) <= dataBufferIn_long(1489);
	dataBufferOut_long(1150) <= dataBufferIn_long(1490);
	dataBufferOut_long(1893) <= dataBufferIn_long(1491);
	dataBufferOut_long(2636) <= dataBufferIn_long(1492);
	dataBufferOut_long(3379) <= dataBufferIn_long(1493);
	dataBufferOut_long(4122) <= dataBufferIn_long(1494);
	dataBufferOut_long(4865) <= dataBufferIn_long(1495);
	dataBufferOut_long(5608) <= dataBufferIn_long(1496);
	dataBufferOut_long( 207) <= dataBufferIn_long(1497);
	dataBufferOut_long( 950) <= dataBufferIn_long(1498);
	dataBufferOut_long(1693) <= dataBufferIn_long(1499);
	dataBufferOut_long(2436) <= dataBufferIn_long(1500);
	dataBufferOut_long(3179) <= dataBufferIn_long(1501);
	dataBufferOut_long(3922) <= dataBufferIn_long(1502);
	dataBufferOut_long(4665) <= dataBufferIn_long(1503);
	dataBufferOut_long(5408) <= dataBufferIn_long(1504);
	dataBufferOut_long(   7) <= dataBufferIn_long(1505);
	dataBufferOut_long( 750) <= dataBufferIn_long(1506);
	dataBufferOut_long(1493) <= dataBufferIn_long(1507);
	dataBufferOut_long(2236) <= dataBufferIn_long(1508);
	dataBufferOut_long(2979) <= dataBufferIn_long(1509);
	dataBufferOut_long(3722) <= dataBufferIn_long(1510);
	dataBufferOut_long(4465) <= dataBufferIn_long(1511);
	dataBufferOut_long(5208) <= dataBufferIn_long(1512);
	dataBufferOut_long(5951) <= dataBufferIn_long(1513);
	dataBufferOut_long( 550) <= dataBufferIn_long(1514);
	dataBufferOut_long(1293) <= dataBufferIn_long(1515);
	dataBufferOut_long(2036) <= dataBufferIn_long(1516);
	dataBufferOut_long(2779) <= dataBufferIn_long(1517);
	dataBufferOut_long(3522) <= dataBufferIn_long(1518);
	dataBufferOut_long(4265) <= dataBufferIn_long(1519);
	dataBufferOut_long(5008) <= dataBufferIn_long(1520);
	dataBufferOut_long(5751) <= dataBufferIn_long(1521);
	dataBufferOut_long( 350) <= dataBufferIn_long(1522);
	dataBufferOut_long(1093) <= dataBufferIn_long(1523);
	dataBufferOut_long(1836) <= dataBufferIn_long(1524);
	dataBufferOut_long(2579) <= dataBufferIn_long(1525);
	dataBufferOut_long(3322) <= dataBufferIn_long(1526);
	dataBufferOut_long(4065) <= dataBufferIn_long(1527);
	dataBufferOut_long(4808) <= dataBufferIn_long(1528);
	dataBufferOut_long(5551) <= dataBufferIn_long(1529);
	dataBufferOut_long( 150) <= dataBufferIn_long(1530);
	dataBufferOut_long( 893) <= dataBufferIn_long(1531);
	dataBufferOut_long(1636) <= dataBufferIn_long(1532);
	dataBufferOut_long(2379) <= dataBufferIn_long(1533);
	dataBufferOut_long(3122) <= dataBufferIn_long(1534);
	dataBufferOut_long(3865) <= dataBufferIn_long(1535);
	dataBufferOut_long(4608) <= dataBufferIn_long(1536);
	dataBufferOut_long(5351) <= dataBufferIn_long(1537);
	dataBufferOut_long(6094) <= dataBufferIn_long(1538);
	dataBufferOut_long( 693) <= dataBufferIn_long(1539);
	dataBufferOut_long(1436) <= dataBufferIn_long(1540);
	dataBufferOut_long(2179) <= dataBufferIn_long(1541);
	dataBufferOut_long(2922) <= dataBufferIn_long(1542);
	dataBufferOut_long(3665) <= dataBufferIn_long(1543);
	dataBufferOut_long(4408) <= dataBufferIn_long(1544);
	dataBufferOut_long(5151) <= dataBufferIn_long(1545);
	dataBufferOut_long(5894) <= dataBufferIn_long(1546);
	dataBufferOut_long( 493) <= dataBufferIn_long(1547);
	dataBufferOut_long(1236) <= dataBufferIn_long(1548);
	dataBufferOut_long(1979) <= dataBufferIn_long(1549);
	dataBufferOut_long(2722) <= dataBufferIn_long(1550);
	dataBufferOut_long(3465) <= dataBufferIn_long(1551);
	dataBufferOut_long(4208) <= dataBufferIn_long(1552);
	dataBufferOut_long(4951) <= dataBufferIn_long(1553);
	dataBufferOut_long(5694) <= dataBufferIn_long(1554);
	dataBufferOut_long( 293) <= dataBufferIn_long(1555);
	dataBufferOut_long(1036) <= dataBufferIn_long(1556);
	dataBufferOut_long(1779) <= dataBufferIn_long(1557);
	dataBufferOut_long(2522) <= dataBufferIn_long(1558);
	dataBufferOut_long(3265) <= dataBufferIn_long(1559);
	dataBufferOut_long(4008) <= dataBufferIn_long(1560);
	dataBufferOut_long(4751) <= dataBufferIn_long(1561);
	dataBufferOut_long(5494) <= dataBufferIn_long(1562);
	dataBufferOut_long(  93) <= dataBufferIn_long(1563);
	dataBufferOut_long( 836) <= dataBufferIn_long(1564);
	dataBufferOut_long(1579) <= dataBufferIn_long(1565);
	dataBufferOut_long(2322) <= dataBufferIn_long(1566);
	dataBufferOut_long(3065) <= dataBufferIn_long(1567);
	dataBufferOut_long(3808) <= dataBufferIn_long(1568);
	dataBufferOut_long(4551) <= dataBufferIn_long(1569);
	dataBufferOut_long(5294) <= dataBufferIn_long(1570);
	dataBufferOut_long(6037) <= dataBufferIn_long(1571);
	dataBufferOut_long( 636) <= dataBufferIn_long(1572);
	dataBufferOut_long(1379) <= dataBufferIn_long(1573);
	dataBufferOut_long(2122) <= dataBufferIn_long(1574);
	dataBufferOut_long(2865) <= dataBufferIn_long(1575);
	dataBufferOut_long(3608) <= dataBufferIn_long(1576);
	dataBufferOut_long(4351) <= dataBufferIn_long(1577);
	dataBufferOut_long(5094) <= dataBufferIn_long(1578);
	dataBufferOut_long(5837) <= dataBufferIn_long(1579);
	dataBufferOut_long( 436) <= dataBufferIn_long(1580);
	dataBufferOut_long(1179) <= dataBufferIn_long(1581);
	dataBufferOut_long(1922) <= dataBufferIn_long(1582);
	dataBufferOut_long(2665) <= dataBufferIn_long(1583);
	dataBufferOut_long(3408) <= dataBufferIn_long(1584);
	dataBufferOut_long(4151) <= dataBufferIn_long(1585);
	dataBufferOut_long(4894) <= dataBufferIn_long(1586);
	dataBufferOut_long(5637) <= dataBufferIn_long(1587);
	dataBufferOut_long( 236) <= dataBufferIn_long(1588);
	dataBufferOut_long( 979) <= dataBufferIn_long(1589);
	dataBufferOut_long(1722) <= dataBufferIn_long(1590);
	dataBufferOut_long(2465) <= dataBufferIn_long(1591);
	dataBufferOut_long(3208) <= dataBufferIn_long(1592);
	dataBufferOut_long(3951) <= dataBufferIn_long(1593);
	dataBufferOut_long(4694) <= dataBufferIn_long(1594);
	dataBufferOut_long(5437) <= dataBufferIn_long(1595);
	dataBufferOut_long(  36) <= dataBufferIn_long(1596);
	dataBufferOut_long( 779) <= dataBufferIn_long(1597);
	dataBufferOut_long(1522) <= dataBufferIn_long(1598);
	dataBufferOut_long(2265) <= dataBufferIn_long(1599);
	dataBufferOut_long(3008) <= dataBufferIn_long(1600);
	dataBufferOut_long(3751) <= dataBufferIn_long(1601);
	dataBufferOut_long(4494) <= dataBufferIn_long(1602);
	dataBufferOut_long(5237) <= dataBufferIn_long(1603);
	dataBufferOut_long(5980) <= dataBufferIn_long(1604);
	dataBufferOut_long( 579) <= dataBufferIn_long(1605);
	dataBufferOut_long(1322) <= dataBufferIn_long(1606);
	dataBufferOut_long(2065) <= dataBufferIn_long(1607);
	dataBufferOut_long(2808) <= dataBufferIn_long(1608);
	dataBufferOut_long(3551) <= dataBufferIn_long(1609);
	dataBufferOut_long(4294) <= dataBufferIn_long(1610);
	dataBufferOut_long(5037) <= dataBufferIn_long(1611);
	dataBufferOut_long(5780) <= dataBufferIn_long(1612);
	dataBufferOut_long( 379) <= dataBufferIn_long(1613);
	dataBufferOut_long(1122) <= dataBufferIn_long(1614);
	dataBufferOut_long(1865) <= dataBufferIn_long(1615);
	dataBufferOut_long(2608) <= dataBufferIn_long(1616);
	dataBufferOut_long(3351) <= dataBufferIn_long(1617);
	dataBufferOut_long(4094) <= dataBufferIn_long(1618);
	dataBufferOut_long(4837) <= dataBufferIn_long(1619);
	dataBufferOut_long(5580) <= dataBufferIn_long(1620);
	dataBufferOut_long( 179) <= dataBufferIn_long(1621);
	dataBufferOut_long( 922) <= dataBufferIn_long(1622);
	dataBufferOut_long(1665) <= dataBufferIn_long(1623);
	dataBufferOut_long(2408) <= dataBufferIn_long(1624);
	dataBufferOut_long(3151) <= dataBufferIn_long(1625);
	dataBufferOut_long(3894) <= dataBufferIn_long(1626);
	dataBufferOut_long(4637) <= dataBufferIn_long(1627);
	dataBufferOut_long(5380) <= dataBufferIn_long(1628);
	dataBufferOut_long(6123) <= dataBufferIn_long(1629);
	dataBufferOut_long( 722) <= dataBufferIn_long(1630);
	dataBufferOut_long(1465) <= dataBufferIn_long(1631);
	dataBufferOut_long(2208) <= dataBufferIn_long(1632);
	dataBufferOut_long(2951) <= dataBufferIn_long(1633);
	dataBufferOut_long(3694) <= dataBufferIn_long(1634);
	dataBufferOut_long(4437) <= dataBufferIn_long(1635);
	dataBufferOut_long(5180) <= dataBufferIn_long(1636);
	dataBufferOut_long(5923) <= dataBufferIn_long(1637);
	dataBufferOut_long( 522) <= dataBufferIn_long(1638);
	dataBufferOut_long(1265) <= dataBufferIn_long(1639);
	dataBufferOut_long(2008) <= dataBufferIn_long(1640);
	dataBufferOut_long(2751) <= dataBufferIn_long(1641);
	dataBufferOut_long(3494) <= dataBufferIn_long(1642);
	dataBufferOut_long(4237) <= dataBufferIn_long(1643);
	dataBufferOut_long(4980) <= dataBufferIn_long(1644);
	dataBufferOut_long(5723) <= dataBufferIn_long(1645);
	dataBufferOut_long( 322) <= dataBufferIn_long(1646);
	dataBufferOut_long(1065) <= dataBufferIn_long(1647);
	dataBufferOut_long(1808) <= dataBufferIn_long(1648);
	dataBufferOut_long(2551) <= dataBufferIn_long(1649);
	dataBufferOut_long(3294) <= dataBufferIn_long(1650);
	dataBufferOut_long(4037) <= dataBufferIn_long(1651);
	dataBufferOut_long(4780) <= dataBufferIn_long(1652);
	dataBufferOut_long(5523) <= dataBufferIn_long(1653);
	dataBufferOut_long( 122) <= dataBufferIn_long(1654);
	dataBufferOut_long( 865) <= dataBufferIn_long(1655);
	dataBufferOut_long(1608) <= dataBufferIn_long(1656);
	dataBufferOut_long(2351) <= dataBufferIn_long(1657);
	dataBufferOut_long(3094) <= dataBufferIn_long(1658);
	dataBufferOut_long(3837) <= dataBufferIn_long(1659);
	dataBufferOut_long(4580) <= dataBufferIn_long(1660);
	dataBufferOut_long(5323) <= dataBufferIn_long(1661);
	dataBufferOut_long(6066) <= dataBufferIn_long(1662);
	dataBufferOut_long( 665) <= dataBufferIn_long(1663);
	dataBufferOut_long(1408) <= dataBufferIn_long(1664);
	dataBufferOut_long(2151) <= dataBufferIn_long(1665);
	dataBufferOut_long(2894) <= dataBufferIn_long(1666);
	dataBufferOut_long(3637) <= dataBufferIn_long(1667);
	dataBufferOut_long(4380) <= dataBufferIn_long(1668);
	dataBufferOut_long(5123) <= dataBufferIn_long(1669);
	dataBufferOut_long(5866) <= dataBufferIn_long(1670);
	dataBufferOut_long( 465) <= dataBufferIn_long(1671);
	dataBufferOut_long(1208) <= dataBufferIn_long(1672);
	dataBufferOut_long(1951) <= dataBufferIn_long(1673);
	dataBufferOut_long(2694) <= dataBufferIn_long(1674);
	dataBufferOut_long(3437) <= dataBufferIn_long(1675);
	dataBufferOut_long(4180) <= dataBufferIn_long(1676);
	dataBufferOut_long(4923) <= dataBufferIn_long(1677);
	dataBufferOut_long(5666) <= dataBufferIn_long(1678);
	dataBufferOut_long( 265) <= dataBufferIn_long(1679);
	dataBufferOut_long(1008) <= dataBufferIn_long(1680);
	dataBufferOut_long(1751) <= dataBufferIn_long(1681);
	dataBufferOut_long(2494) <= dataBufferIn_long(1682);
	dataBufferOut_long(3237) <= dataBufferIn_long(1683);
	dataBufferOut_long(3980) <= dataBufferIn_long(1684);
	dataBufferOut_long(4723) <= dataBufferIn_long(1685);
	dataBufferOut_long(5466) <= dataBufferIn_long(1686);
	dataBufferOut_long(  65) <= dataBufferIn_long(1687);
	dataBufferOut_long( 808) <= dataBufferIn_long(1688);
	dataBufferOut_long(1551) <= dataBufferIn_long(1689);
	dataBufferOut_long(2294) <= dataBufferIn_long(1690);
	dataBufferOut_long(3037) <= dataBufferIn_long(1691);
	dataBufferOut_long(3780) <= dataBufferIn_long(1692);
	dataBufferOut_long(4523) <= dataBufferIn_long(1693);
	dataBufferOut_long(5266) <= dataBufferIn_long(1694);
	dataBufferOut_long(6009) <= dataBufferIn_long(1695);
	dataBufferOut_long( 608) <= dataBufferIn_long(1696);
	dataBufferOut_long(1351) <= dataBufferIn_long(1697);
	dataBufferOut_long(2094) <= dataBufferIn_long(1698);
	dataBufferOut_long(2837) <= dataBufferIn_long(1699);
	dataBufferOut_long(3580) <= dataBufferIn_long(1700);
	dataBufferOut_long(4323) <= dataBufferIn_long(1701);
	dataBufferOut_long(5066) <= dataBufferIn_long(1702);
	dataBufferOut_long(5809) <= dataBufferIn_long(1703);
	dataBufferOut_long( 408) <= dataBufferIn_long(1704);
	dataBufferOut_long(1151) <= dataBufferIn_long(1705);
	dataBufferOut_long(1894) <= dataBufferIn_long(1706);
	dataBufferOut_long(2637) <= dataBufferIn_long(1707);
	dataBufferOut_long(3380) <= dataBufferIn_long(1708);
	dataBufferOut_long(4123) <= dataBufferIn_long(1709);
	dataBufferOut_long(4866) <= dataBufferIn_long(1710);
	dataBufferOut_long(5609) <= dataBufferIn_long(1711);
	dataBufferOut_long( 208) <= dataBufferIn_long(1712);
	dataBufferOut_long( 951) <= dataBufferIn_long(1713);
	dataBufferOut_long(1694) <= dataBufferIn_long(1714);
	dataBufferOut_long(2437) <= dataBufferIn_long(1715);
	dataBufferOut_long(3180) <= dataBufferIn_long(1716);
	dataBufferOut_long(3923) <= dataBufferIn_long(1717);
	dataBufferOut_long(4666) <= dataBufferIn_long(1718);
	dataBufferOut_long(5409) <= dataBufferIn_long(1719);
	dataBufferOut_long(   8) <= dataBufferIn_long(1720);
	dataBufferOut_long( 751) <= dataBufferIn_long(1721);
	dataBufferOut_long(1494) <= dataBufferIn_long(1722);
	dataBufferOut_long(2237) <= dataBufferIn_long(1723);
	dataBufferOut_long(2980) <= dataBufferIn_long(1724);
	dataBufferOut_long(3723) <= dataBufferIn_long(1725);
	dataBufferOut_long(4466) <= dataBufferIn_long(1726);
	dataBufferOut_long(5209) <= dataBufferIn_long(1727);
	dataBufferOut_long(5952) <= dataBufferIn_long(1728);
	dataBufferOut_long( 551) <= dataBufferIn_long(1729);
	dataBufferOut_long(1294) <= dataBufferIn_long(1730);
	dataBufferOut_long(2037) <= dataBufferIn_long(1731);
	dataBufferOut_long(2780) <= dataBufferIn_long(1732);
	dataBufferOut_long(3523) <= dataBufferIn_long(1733);
	dataBufferOut_long(4266) <= dataBufferIn_long(1734);
	dataBufferOut_long(5009) <= dataBufferIn_long(1735);
	dataBufferOut_long(5752) <= dataBufferIn_long(1736);
	dataBufferOut_long( 351) <= dataBufferIn_long(1737);
	dataBufferOut_long(1094) <= dataBufferIn_long(1738);
	dataBufferOut_long(1837) <= dataBufferIn_long(1739);
	dataBufferOut_long(2580) <= dataBufferIn_long(1740);
	dataBufferOut_long(3323) <= dataBufferIn_long(1741);
	dataBufferOut_long(4066) <= dataBufferIn_long(1742);
	dataBufferOut_long(4809) <= dataBufferIn_long(1743);
	dataBufferOut_long(5552) <= dataBufferIn_long(1744);
	dataBufferOut_long( 151) <= dataBufferIn_long(1745);
	dataBufferOut_long( 894) <= dataBufferIn_long(1746);
	dataBufferOut_long(1637) <= dataBufferIn_long(1747);
	dataBufferOut_long(2380) <= dataBufferIn_long(1748);
	dataBufferOut_long(3123) <= dataBufferIn_long(1749);
	dataBufferOut_long(3866) <= dataBufferIn_long(1750);
	dataBufferOut_long(4609) <= dataBufferIn_long(1751);
	dataBufferOut_long(5352) <= dataBufferIn_long(1752);
	dataBufferOut_long(6095) <= dataBufferIn_long(1753);
	dataBufferOut_long( 694) <= dataBufferIn_long(1754);
	dataBufferOut_long(1437) <= dataBufferIn_long(1755);
	dataBufferOut_long(2180) <= dataBufferIn_long(1756);
	dataBufferOut_long(2923) <= dataBufferIn_long(1757);
	dataBufferOut_long(3666) <= dataBufferIn_long(1758);
	dataBufferOut_long(4409) <= dataBufferIn_long(1759);
	dataBufferOut_long(5152) <= dataBufferIn_long(1760);
	dataBufferOut_long(5895) <= dataBufferIn_long(1761);
	dataBufferOut_long( 494) <= dataBufferIn_long(1762);
	dataBufferOut_long(1237) <= dataBufferIn_long(1763);
	dataBufferOut_long(1980) <= dataBufferIn_long(1764);
	dataBufferOut_long(2723) <= dataBufferIn_long(1765);
	dataBufferOut_long(3466) <= dataBufferIn_long(1766);
	dataBufferOut_long(4209) <= dataBufferIn_long(1767);
	dataBufferOut_long(4952) <= dataBufferIn_long(1768);
	dataBufferOut_long(5695) <= dataBufferIn_long(1769);
	dataBufferOut_long( 294) <= dataBufferIn_long(1770);
	dataBufferOut_long(1037) <= dataBufferIn_long(1771);
	dataBufferOut_long(1780) <= dataBufferIn_long(1772);
	dataBufferOut_long(2523) <= dataBufferIn_long(1773);
	dataBufferOut_long(3266) <= dataBufferIn_long(1774);
	dataBufferOut_long(4009) <= dataBufferIn_long(1775);
	dataBufferOut_long(4752) <= dataBufferIn_long(1776);
	dataBufferOut_long(5495) <= dataBufferIn_long(1777);
	dataBufferOut_long(  94) <= dataBufferIn_long(1778);
	dataBufferOut_long( 837) <= dataBufferIn_long(1779);
	dataBufferOut_long(1580) <= dataBufferIn_long(1780);
	dataBufferOut_long(2323) <= dataBufferIn_long(1781);
	dataBufferOut_long(3066) <= dataBufferIn_long(1782);
	dataBufferOut_long(3809) <= dataBufferIn_long(1783);
	dataBufferOut_long(4552) <= dataBufferIn_long(1784);
	dataBufferOut_long(5295) <= dataBufferIn_long(1785);
	dataBufferOut_long(6038) <= dataBufferIn_long(1786);
	dataBufferOut_long( 637) <= dataBufferIn_long(1787);
	dataBufferOut_long(1380) <= dataBufferIn_long(1788);
	dataBufferOut_long(2123) <= dataBufferIn_long(1789);
	dataBufferOut_long(2866) <= dataBufferIn_long(1790);
	dataBufferOut_long(3609) <= dataBufferIn_long(1791);
	dataBufferOut_long(4352) <= dataBufferIn_long(1792);
	dataBufferOut_long(5095) <= dataBufferIn_long(1793);
	dataBufferOut_long(5838) <= dataBufferIn_long(1794);
	dataBufferOut_long( 437) <= dataBufferIn_long(1795);
	dataBufferOut_long(1180) <= dataBufferIn_long(1796);
	dataBufferOut_long(1923) <= dataBufferIn_long(1797);
	dataBufferOut_long(2666) <= dataBufferIn_long(1798);
	dataBufferOut_long(3409) <= dataBufferIn_long(1799);
	dataBufferOut_long(4152) <= dataBufferIn_long(1800);
	dataBufferOut_long(4895) <= dataBufferIn_long(1801);
	dataBufferOut_long(5638) <= dataBufferIn_long(1802);
	dataBufferOut_long( 237) <= dataBufferIn_long(1803);
	dataBufferOut_long( 980) <= dataBufferIn_long(1804);
	dataBufferOut_long(1723) <= dataBufferIn_long(1805);
	dataBufferOut_long(2466) <= dataBufferIn_long(1806);
	dataBufferOut_long(3209) <= dataBufferIn_long(1807);
	dataBufferOut_long(3952) <= dataBufferIn_long(1808);
	dataBufferOut_long(4695) <= dataBufferIn_long(1809);
	dataBufferOut_long(5438) <= dataBufferIn_long(1810);
	dataBufferOut_long(  37) <= dataBufferIn_long(1811);
	dataBufferOut_long( 780) <= dataBufferIn_long(1812);
	dataBufferOut_long(1523) <= dataBufferIn_long(1813);
	dataBufferOut_long(2266) <= dataBufferIn_long(1814);
	dataBufferOut_long(3009) <= dataBufferIn_long(1815);
	dataBufferOut_long(3752) <= dataBufferIn_long(1816);
	dataBufferOut_long(4495) <= dataBufferIn_long(1817);
	dataBufferOut_long(5238) <= dataBufferIn_long(1818);
	dataBufferOut_long(5981) <= dataBufferIn_long(1819);
	dataBufferOut_long( 580) <= dataBufferIn_long(1820);
	dataBufferOut_long(1323) <= dataBufferIn_long(1821);
	dataBufferOut_long(2066) <= dataBufferIn_long(1822);
	dataBufferOut_long(2809) <= dataBufferIn_long(1823);
	dataBufferOut_long(3552) <= dataBufferIn_long(1824);
	dataBufferOut_long(4295) <= dataBufferIn_long(1825);
	dataBufferOut_long(5038) <= dataBufferIn_long(1826);
	dataBufferOut_long(5781) <= dataBufferIn_long(1827);
	dataBufferOut_long( 380) <= dataBufferIn_long(1828);
	dataBufferOut_long(1123) <= dataBufferIn_long(1829);
	dataBufferOut_long(1866) <= dataBufferIn_long(1830);
	dataBufferOut_long(2609) <= dataBufferIn_long(1831);
	dataBufferOut_long(3352) <= dataBufferIn_long(1832);
	dataBufferOut_long(4095) <= dataBufferIn_long(1833);
	dataBufferOut_long(4838) <= dataBufferIn_long(1834);
	dataBufferOut_long(5581) <= dataBufferIn_long(1835);
	dataBufferOut_long( 180) <= dataBufferIn_long(1836);
	dataBufferOut_long( 923) <= dataBufferIn_long(1837);
	dataBufferOut_long(1666) <= dataBufferIn_long(1838);
	dataBufferOut_long(2409) <= dataBufferIn_long(1839);
	dataBufferOut_long(3152) <= dataBufferIn_long(1840);
	dataBufferOut_long(3895) <= dataBufferIn_long(1841);
	dataBufferOut_long(4638) <= dataBufferIn_long(1842);
	dataBufferOut_long(5381) <= dataBufferIn_long(1843);
	dataBufferOut_long(6124) <= dataBufferIn_long(1844);
	dataBufferOut_long( 723) <= dataBufferIn_long(1845);
	dataBufferOut_long(1466) <= dataBufferIn_long(1846);
	dataBufferOut_long(2209) <= dataBufferIn_long(1847);
	dataBufferOut_long(2952) <= dataBufferIn_long(1848);
	dataBufferOut_long(3695) <= dataBufferIn_long(1849);
	dataBufferOut_long(4438) <= dataBufferIn_long(1850);
	dataBufferOut_long(5181) <= dataBufferIn_long(1851);
	dataBufferOut_long(5924) <= dataBufferIn_long(1852);
	dataBufferOut_long( 523) <= dataBufferIn_long(1853);
	dataBufferOut_long(1266) <= dataBufferIn_long(1854);
	dataBufferOut_long(2009) <= dataBufferIn_long(1855);
	dataBufferOut_long(2752) <= dataBufferIn_long(1856);
	dataBufferOut_long(3495) <= dataBufferIn_long(1857);
	dataBufferOut_long(4238) <= dataBufferIn_long(1858);
	dataBufferOut_long(4981) <= dataBufferIn_long(1859);
	dataBufferOut_long(5724) <= dataBufferIn_long(1860);
	dataBufferOut_long( 323) <= dataBufferIn_long(1861);
	dataBufferOut_long(1066) <= dataBufferIn_long(1862);
	dataBufferOut_long(1809) <= dataBufferIn_long(1863);
	dataBufferOut_long(2552) <= dataBufferIn_long(1864);
	dataBufferOut_long(3295) <= dataBufferIn_long(1865);
	dataBufferOut_long(4038) <= dataBufferIn_long(1866);
	dataBufferOut_long(4781) <= dataBufferIn_long(1867);
	dataBufferOut_long(5524) <= dataBufferIn_long(1868);
	dataBufferOut_long( 123) <= dataBufferIn_long(1869);
	dataBufferOut_long( 866) <= dataBufferIn_long(1870);
	dataBufferOut_long(1609) <= dataBufferIn_long(1871);
	dataBufferOut_long(2352) <= dataBufferIn_long(1872);
	dataBufferOut_long(3095) <= dataBufferIn_long(1873);
	dataBufferOut_long(3838) <= dataBufferIn_long(1874);
	dataBufferOut_long(4581) <= dataBufferIn_long(1875);
	dataBufferOut_long(5324) <= dataBufferIn_long(1876);
	dataBufferOut_long(6067) <= dataBufferIn_long(1877);
	dataBufferOut_long( 666) <= dataBufferIn_long(1878);
	dataBufferOut_long(1409) <= dataBufferIn_long(1879);
	dataBufferOut_long(2152) <= dataBufferIn_long(1880);
	dataBufferOut_long(2895) <= dataBufferIn_long(1881);
	dataBufferOut_long(3638) <= dataBufferIn_long(1882);
	dataBufferOut_long(4381) <= dataBufferIn_long(1883);
	dataBufferOut_long(5124) <= dataBufferIn_long(1884);
	dataBufferOut_long(5867) <= dataBufferIn_long(1885);
	dataBufferOut_long( 466) <= dataBufferIn_long(1886);
	dataBufferOut_long(1209) <= dataBufferIn_long(1887);
	dataBufferOut_long(1952) <= dataBufferIn_long(1888);
	dataBufferOut_long(2695) <= dataBufferIn_long(1889);
	dataBufferOut_long(3438) <= dataBufferIn_long(1890);
	dataBufferOut_long(4181) <= dataBufferIn_long(1891);
	dataBufferOut_long(4924) <= dataBufferIn_long(1892);
	dataBufferOut_long(5667) <= dataBufferIn_long(1893);
	dataBufferOut_long( 266) <= dataBufferIn_long(1894);
	dataBufferOut_long(1009) <= dataBufferIn_long(1895);
	dataBufferOut_long(1752) <= dataBufferIn_long(1896);
	dataBufferOut_long(2495) <= dataBufferIn_long(1897);
	dataBufferOut_long(3238) <= dataBufferIn_long(1898);
	dataBufferOut_long(3981) <= dataBufferIn_long(1899);
	dataBufferOut_long(4724) <= dataBufferIn_long(1900);
	dataBufferOut_long(5467) <= dataBufferIn_long(1901);
	dataBufferOut_long(  66) <= dataBufferIn_long(1902);
	dataBufferOut_long( 809) <= dataBufferIn_long(1903);
	dataBufferOut_long(1552) <= dataBufferIn_long(1904);
	dataBufferOut_long(2295) <= dataBufferIn_long(1905);
	dataBufferOut_long(3038) <= dataBufferIn_long(1906);
	dataBufferOut_long(3781) <= dataBufferIn_long(1907);
	dataBufferOut_long(4524) <= dataBufferIn_long(1908);
	dataBufferOut_long(5267) <= dataBufferIn_long(1909);
	dataBufferOut_long(6010) <= dataBufferIn_long(1910);
	dataBufferOut_long( 609) <= dataBufferIn_long(1911);
	dataBufferOut_long(1352) <= dataBufferIn_long(1912);
	dataBufferOut_long(2095) <= dataBufferIn_long(1913);
	dataBufferOut_long(2838) <= dataBufferIn_long(1914);
	dataBufferOut_long(3581) <= dataBufferIn_long(1915);
	dataBufferOut_long(4324) <= dataBufferIn_long(1916);
	dataBufferOut_long(5067) <= dataBufferIn_long(1917);
	dataBufferOut_long(5810) <= dataBufferIn_long(1918);
	dataBufferOut_long( 409) <= dataBufferIn_long(1919);
	dataBufferOut_long(1152) <= dataBufferIn_long(1920);
	dataBufferOut_long(1895) <= dataBufferIn_long(1921);
	dataBufferOut_long(2638) <= dataBufferIn_long(1922);
	dataBufferOut_long(3381) <= dataBufferIn_long(1923);
	dataBufferOut_long(4124) <= dataBufferIn_long(1924);
	dataBufferOut_long(4867) <= dataBufferIn_long(1925);
	dataBufferOut_long(5610) <= dataBufferIn_long(1926);
	dataBufferOut_long( 209) <= dataBufferIn_long(1927);
	dataBufferOut_long( 952) <= dataBufferIn_long(1928);
	dataBufferOut_long(1695) <= dataBufferIn_long(1929);
	dataBufferOut_long(2438) <= dataBufferIn_long(1930);
	dataBufferOut_long(3181) <= dataBufferIn_long(1931);
	dataBufferOut_long(3924) <= dataBufferIn_long(1932);
	dataBufferOut_long(4667) <= dataBufferIn_long(1933);
	dataBufferOut_long(5410) <= dataBufferIn_long(1934);
	dataBufferOut_long(   9) <= dataBufferIn_long(1935);
	dataBufferOut_long( 752) <= dataBufferIn_long(1936);
	dataBufferOut_long(1495) <= dataBufferIn_long(1937);
	dataBufferOut_long(2238) <= dataBufferIn_long(1938);
	dataBufferOut_long(2981) <= dataBufferIn_long(1939);
	dataBufferOut_long(3724) <= dataBufferIn_long(1940);
	dataBufferOut_long(4467) <= dataBufferIn_long(1941);
	dataBufferOut_long(5210) <= dataBufferIn_long(1942);
	dataBufferOut_long(5953) <= dataBufferIn_long(1943);
	dataBufferOut_long( 552) <= dataBufferIn_long(1944);
	dataBufferOut_long(1295) <= dataBufferIn_long(1945);
	dataBufferOut_long(2038) <= dataBufferIn_long(1946);
	dataBufferOut_long(2781) <= dataBufferIn_long(1947);
	dataBufferOut_long(3524) <= dataBufferIn_long(1948);
	dataBufferOut_long(4267) <= dataBufferIn_long(1949);
	dataBufferOut_long(5010) <= dataBufferIn_long(1950);
	dataBufferOut_long(5753) <= dataBufferIn_long(1951);
	dataBufferOut_long( 352) <= dataBufferIn_long(1952);
	dataBufferOut_long(1095) <= dataBufferIn_long(1953);
	dataBufferOut_long(1838) <= dataBufferIn_long(1954);
	dataBufferOut_long(2581) <= dataBufferIn_long(1955);
	dataBufferOut_long(3324) <= dataBufferIn_long(1956);
	dataBufferOut_long(4067) <= dataBufferIn_long(1957);
	dataBufferOut_long(4810) <= dataBufferIn_long(1958);
	dataBufferOut_long(5553) <= dataBufferIn_long(1959);
	dataBufferOut_long( 152) <= dataBufferIn_long(1960);
	dataBufferOut_long( 895) <= dataBufferIn_long(1961);
	dataBufferOut_long(1638) <= dataBufferIn_long(1962);
	dataBufferOut_long(2381) <= dataBufferIn_long(1963);
	dataBufferOut_long(3124) <= dataBufferIn_long(1964);
	dataBufferOut_long(3867) <= dataBufferIn_long(1965);
	dataBufferOut_long(4610) <= dataBufferIn_long(1966);
	dataBufferOut_long(5353) <= dataBufferIn_long(1967);
	dataBufferOut_long(6096) <= dataBufferIn_long(1968);
	dataBufferOut_long( 695) <= dataBufferIn_long(1969);
	dataBufferOut_long(1438) <= dataBufferIn_long(1970);
	dataBufferOut_long(2181) <= dataBufferIn_long(1971);
	dataBufferOut_long(2924) <= dataBufferIn_long(1972);
	dataBufferOut_long(3667) <= dataBufferIn_long(1973);
	dataBufferOut_long(4410) <= dataBufferIn_long(1974);
	dataBufferOut_long(5153) <= dataBufferIn_long(1975);
	dataBufferOut_long(5896) <= dataBufferIn_long(1976);
	dataBufferOut_long( 495) <= dataBufferIn_long(1977);
	dataBufferOut_long(1238) <= dataBufferIn_long(1978);
	dataBufferOut_long(1981) <= dataBufferIn_long(1979);
	dataBufferOut_long(2724) <= dataBufferIn_long(1980);
	dataBufferOut_long(3467) <= dataBufferIn_long(1981);
	dataBufferOut_long(4210) <= dataBufferIn_long(1982);
	dataBufferOut_long(4953) <= dataBufferIn_long(1983);
	dataBufferOut_long(5696) <= dataBufferIn_long(1984);
	dataBufferOut_long( 295) <= dataBufferIn_long(1985);
	dataBufferOut_long(1038) <= dataBufferIn_long(1986);
	dataBufferOut_long(1781) <= dataBufferIn_long(1987);
	dataBufferOut_long(2524) <= dataBufferIn_long(1988);
	dataBufferOut_long(3267) <= dataBufferIn_long(1989);
	dataBufferOut_long(4010) <= dataBufferIn_long(1990);
	dataBufferOut_long(4753) <= dataBufferIn_long(1991);
	dataBufferOut_long(5496) <= dataBufferIn_long(1992);
	dataBufferOut_long(  95) <= dataBufferIn_long(1993);
	dataBufferOut_long( 838) <= dataBufferIn_long(1994);
	dataBufferOut_long(1581) <= dataBufferIn_long(1995);
	dataBufferOut_long(2324) <= dataBufferIn_long(1996);
	dataBufferOut_long(3067) <= dataBufferIn_long(1997);
	dataBufferOut_long(3810) <= dataBufferIn_long(1998);
	dataBufferOut_long(4553) <= dataBufferIn_long(1999);
	dataBufferOut_long(5296) <= dataBufferIn_long(2000);
	dataBufferOut_long(6039) <= dataBufferIn_long(2001);
	dataBufferOut_long( 638) <= dataBufferIn_long(2002);
	dataBufferOut_long(1381) <= dataBufferIn_long(2003);
	dataBufferOut_long(2124) <= dataBufferIn_long(2004);
	dataBufferOut_long(2867) <= dataBufferIn_long(2005);
	dataBufferOut_long(3610) <= dataBufferIn_long(2006);
	dataBufferOut_long(4353) <= dataBufferIn_long(2007);
	dataBufferOut_long(5096) <= dataBufferIn_long(2008);
	dataBufferOut_long(5839) <= dataBufferIn_long(2009);
	dataBufferOut_long( 438) <= dataBufferIn_long(2010);
	dataBufferOut_long(1181) <= dataBufferIn_long(2011);
	dataBufferOut_long(1924) <= dataBufferIn_long(2012);
	dataBufferOut_long(2667) <= dataBufferIn_long(2013);
	dataBufferOut_long(3410) <= dataBufferIn_long(2014);
	dataBufferOut_long(4153) <= dataBufferIn_long(2015);
	dataBufferOut_long(4896) <= dataBufferIn_long(2016);
	dataBufferOut_long(5639) <= dataBufferIn_long(2017);
	dataBufferOut_long( 238) <= dataBufferIn_long(2018);
	dataBufferOut_long( 981) <= dataBufferIn_long(2019);
	dataBufferOut_long(1724) <= dataBufferIn_long(2020);
	dataBufferOut_long(2467) <= dataBufferIn_long(2021);
	dataBufferOut_long(3210) <= dataBufferIn_long(2022);
	dataBufferOut_long(3953) <= dataBufferIn_long(2023);
	dataBufferOut_long(4696) <= dataBufferIn_long(2024);
	dataBufferOut_long(5439) <= dataBufferIn_long(2025);
	dataBufferOut_long(  38) <= dataBufferIn_long(2026);
	dataBufferOut_long( 781) <= dataBufferIn_long(2027);
	dataBufferOut_long(1524) <= dataBufferIn_long(2028);
	dataBufferOut_long(2267) <= dataBufferIn_long(2029);
	dataBufferOut_long(3010) <= dataBufferIn_long(2030);
	dataBufferOut_long(3753) <= dataBufferIn_long(2031);
	dataBufferOut_long(4496) <= dataBufferIn_long(2032);
	dataBufferOut_long(5239) <= dataBufferIn_long(2033);
	dataBufferOut_long(5982) <= dataBufferIn_long(2034);
	dataBufferOut_long( 581) <= dataBufferIn_long(2035);
	dataBufferOut_long(1324) <= dataBufferIn_long(2036);
	dataBufferOut_long(2067) <= dataBufferIn_long(2037);
	dataBufferOut_long(2810) <= dataBufferIn_long(2038);
	dataBufferOut_long(3553) <= dataBufferIn_long(2039);
	dataBufferOut_long(4296) <= dataBufferIn_long(2040);
	dataBufferOut_long(5039) <= dataBufferIn_long(2041);
	dataBufferOut_long(5782) <= dataBufferIn_long(2042);
	dataBufferOut_long( 381) <= dataBufferIn_long(2043);
	dataBufferOut_long(1124) <= dataBufferIn_long(2044);
	dataBufferOut_long(1867) <= dataBufferIn_long(2045);
	dataBufferOut_long(2610) <= dataBufferIn_long(2046);
	dataBufferOut_long(3353) <= dataBufferIn_long(2047);
	dataBufferOut_long(4096) <= dataBufferIn_long(2048);
	dataBufferOut_long(4839) <= dataBufferIn_long(2049);
	dataBufferOut_long(5582) <= dataBufferIn_long(2050);
	dataBufferOut_long( 181) <= dataBufferIn_long(2051);
	dataBufferOut_long( 924) <= dataBufferIn_long(2052);
	dataBufferOut_long(1667) <= dataBufferIn_long(2053);
	dataBufferOut_long(2410) <= dataBufferIn_long(2054);
	dataBufferOut_long(3153) <= dataBufferIn_long(2055);
	dataBufferOut_long(3896) <= dataBufferIn_long(2056);
	dataBufferOut_long(4639) <= dataBufferIn_long(2057);
	dataBufferOut_long(5382) <= dataBufferIn_long(2058);
	dataBufferOut_long(6125) <= dataBufferIn_long(2059);
	dataBufferOut_long( 724) <= dataBufferIn_long(2060);
	dataBufferOut_long(1467) <= dataBufferIn_long(2061);
	dataBufferOut_long(2210) <= dataBufferIn_long(2062);
	dataBufferOut_long(2953) <= dataBufferIn_long(2063);
	dataBufferOut_long(3696) <= dataBufferIn_long(2064);
	dataBufferOut_long(4439) <= dataBufferIn_long(2065);
	dataBufferOut_long(5182) <= dataBufferIn_long(2066);
	dataBufferOut_long(5925) <= dataBufferIn_long(2067);
	dataBufferOut_long( 524) <= dataBufferIn_long(2068);
	dataBufferOut_long(1267) <= dataBufferIn_long(2069);
	dataBufferOut_long(2010) <= dataBufferIn_long(2070);
	dataBufferOut_long(2753) <= dataBufferIn_long(2071);
	dataBufferOut_long(3496) <= dataBufferIn_long(2072);
	dataBufferOut_long(4239) <= dataBufferIn_long(2073);
	dataBufferOut_long(4982) <= dataBufferIn_long(2074);
	dataBufferOut_long(5725) <= dataBufferIn_long(2075);
	dataBufferOut_long( 324) <= dataBufferIn_long(2076);
	dataBufferOut_long(1067) <= dataBufferIn_long(2077);
	dataBufferOut_long(1810) <= dataBufferIn_long(2078);
	dataBufferOut_long(2553) <= dataBufferIn_long(2079);
	dataBufferOut_long(3296) <= dataBufferIn_long(2080);
	dataBufferOut_long(4039) <= dataBufferIn_long(2081);
	dataBufferOut_long(4782) <= dataBufferIn_long(2082);
	dataBufferOut_long(5525) <= dataBufferIn_long(2083);
	dataBufferOut_long( 124) <= dataBufferIn_long(2084);
	dataBufferOut_long( 867) <= dataBufferIn_long(2085);
	dataBufferOut_long(1610) <= dataBufferIn_long(2086);
	dataBufferOut_long(2353) <= dataBufferIn_long(2087);
	dataBufferOut_long(3096) <= dataBufferIn_long(2088);
	dataBufferOut_long(3839) <= dataBufferIn_long(2089);
	dataBufferOut_long(4582) <= dataBufferIn_long(2090);
	dataBufferOut_long(5325) <= dataBufferIn_long(2091);
	dataBufferOut_long(6068) <= dataBufferIn_long(2092);
	dataBufferOut_long( 667) <= dataBufferIn_long(2093);
	dataBufferOut_long(1410) <= dataBufferIn_long(2094);
	dataBufferOut_long(2153) <= dataBufferIn_long(2095);
	dataBufferOut_long(2896) <= dataBufferIn_long(2096);
	dataBufferOut_long(3639) <= dataBufferIn_long(2097);
	dataBufferOut_long(4382) <= dataBufferIn_long(2098);
	dataBufferOut_long(5125) <= dataBufferIn_long(2099);
	dataBufferOut_long(5868) <= dataBufferIn_long(2100);
	dataBufferOut_long( 467) <= dataBufferIn_long(2101);
	dataBufferOut_long(1210) <= dataBufferIn_long(2102);
	dataBufferOut_long(1953) <= dataBufferIn_long(2103);
	dataBufferOut_long(2696) <= dataBufferIn_long(2104);
	dataBufferOut_long(3439) <= dataBufferIn_long(2105);
	dataBufferOut_long(4182) <= dataBufferIn_long(2106);
	dataBufferOut_long(4925) <= dataBufferIn_long(2107);
	dataBufferOut_long(5668) <= dataBufferIn_long(2108);
	dataBufferOut_long( 267) <= dataBufferIn_long(2109);
	dataBufferOut_long(1010) <= dataBufferIn_long(2110);
	dataBufferOut_long(1753) <= dataBufferIn_long(2111);
	dataBufferOut_long(2496) <= dataBufferIn_long(2112);
	dataBufferOut_long(3239) <= dataBufferIn_long(2113);
	dataBufferOut_long(3982) <= dataBufferIn_long(2114);
	dataBufferOut_long(4725) <= dataBufferIn_long(2115);
	dataBufferOut_long(5468) <= dataBufferIn_long(2116);
	dataBufferOut_long(  67) <= dataBufferIn_long(2117);
	dataBufferOut_long( 810) <= dataBufferIn_long(2118);
	dataBufferOut_long(1553) <= dataBufferIn_long(2119);
	dataBufferOut_long(2296) <= dataBufferIn_long(2120);
	dataBufferOut_long(3039) <= dataBufferIn_long(2121);
	dataBufferOut_long(3782) <= dataBufferIn_long(2122);
	dataBufferOut_long(4525) <= dataBufferIn_long(2123);
	dataBufferOut_long(5268) <= dataBufferIn_long(2124);
	dataBufferOut_long(6011) <= dataBufferIn_long(2125);
	dataBufferOut_long( 610) <= dataBufferIn_long(2126);
	dataBufferOut_long(1353) <= dataBufferIn_long(2127);
	dataBufferOut_long(2096) <= dataBufferIn_long(2128);
	dataBufferOut_long(2839) <= dataBufferIn_long(2129);
	dataBufferOut_long(3582) <= dataBufferIn_long(2130);
	dataBufferOut_long(4325) <= dataBufferIn_long(2131);
	dataBufferOut_long(5068) <= dataBufferIn_long(2132);
	dataBufferOut_long(5811) <= dataBufferIn_long(2133);
	dataBufferOut_long( 410) <= dataBufferIn_long(2134);
	dataBufferOut_long(1153) <= dataBufferIn_long(2135);
	dataBufferOut_long(1896) <= dataBufferIn_long(2136);
	dataBufferOut_long(2639) <= dataBufferIn_long(2137);
	dataBufferOut_long(3382) <= dataBufferIn_long(2138);
	dataBufferOut_long(4125) <= dataBufferIn_long(2139);
	dataBufferOut_long(4868) <= dataBufferIn_long(2140);
	dataBufferOut_long(5611) <= dataBufferIn_long(2141);
	dataBufferOut_long( 210) <= dataBufferIn_long(2142);
	dataBufferOut_long( 953) <= dataBufferIn_long(2143);
	dataBufferOut_long(1696) <= dataBufferIn_long(2144);
	dataBufferOut_long(2439) <= dataBufferIn_long(2145);
	dataBufferOut_long(3182) <= dataBufferIn_long(2146);
	dataBufferOut_long(3925) <= dataBufferIn_long(2147);
	dataBufferOut_long(4668) <= dataBufferIn_long(2148);
	dataBufferOut_long(5411) <= dataBufferIn_long(2149);
	dataBufferOut_long(  10) <= dataBufferIn_long(2150);
	dataBufferOut_long( 753) <= dataBufferIn_long(2151);
	dataBufferOut_long(1496) <= dataBufferIn_long(2152);
	dataBufferOut_long(2239) <= dataBufferIn_long(2153);
	dataBufferOut_long(2982) <= dataBufferIn_long(2154);
	dataBufferOut_long(3725) <= dataBufferIn_long(2155);
	dataBufferOut_long(4468) <= dataBufferIn_long(2156);
	dataBufferOut_long(5211) <= dataBufferIn_long(2157);
	dataBufferOut_long(5954) <= dataBufferIn_long(2158);
	dataBufferOut_long( 553) <= dataBufferIn_long(2159);
	dataBufferOut_long(1296) <= dataBufferIn_long(2160);
	dataBufferOut_long(2039) <= dataBufferIn_long(2161);
	dataBufferOut_long(2782) <= dataBufferIn_long(2162);
	dataBufferOut_long(3525) <= dataBufferIn_long(2163);
	dataBufferOut_long(4268) <= dataBufferIn_long(2164);
	dataBufferOut_long(5011) <= dataBufferIn_long(2165);
	dataBufferOut_long(5754) <= dataBufferIn_long(2166);
	dataBufferOut_long( 353) <= dataBufferIn_long(2167);
	dataBufferOut_long(1096) <= dataBufferIn_long(2168);
	dataBufferOut_long(1839) <= dataBufferIn_long(2169);
	dataBufferOut_long(2582) <= dataBufferIn_long(2170);
	dataBufferOut_long(3325) <= dataBufferIn_long(2171);
	dataBufferOut_long(4068) <= dataBufferIn_long(2172);
	dataBufferOut_long(4811) <= dataBufferIn_long(2173);
	dataBufferOut_long(5554) <= dataBufferIn_long(2174);
	dataBufferOut_long( 153) <= dataBufferIn_long(2175);
	dataBufferOut_long( 896) <= dataBufferIn_long(2176);
	dataBufferOut_long(1639) <= dataBufferIn_long(2177);
	dataBufferOut_long(2382) <= dataBufferIn_long(2178);
	dataBufferOut_long(3125) <= dataBufferIn_long(2179);
	dataBufferOut_long(3868) <= dataBufferIn_long(2180);
	dataBufferOut_long(4611) <= dataBufferIn_long(2181);
	dataBufferOut_long(5354) <= dataBufferIn_long(2182);
	dataBufferOut_long(6097) <= dataBufferIn_long(2183);
	dataBufferOut_long( 696) <= dataBufferIn_long(2184);
	dataBufferOut_long(1439) <= dataBufferIn_long(2185);
	dataBufferOut_long(2182) <= dataBufferIn_long(2186);
	dataBufferOut_long(2925) <= dataBufferIn_long(2187);
	dataBufferOut_long(3668) <= dataBufferIn_long(2188);
	dataBufferOut_long(4411) <= dataBufferIn_long(2189);
	dataBufferOut_long(5154) <= dataBufferIn_long(2190);
	dataBufferOut_long(5897) <= dataBufferIn_long(2191);
	dataBufferOut_long( 496) <= dataBufferIn_long(2192);
	dataBufferOut_long(1239) <= dataBufferIn_long(2193);
	dataBufferOut_long(1982) <= dataBufferIn_long(2194);
	dataBufferOut_long(2725) <= dataBufferIn_long(2195);
	dataBufferOut_long(3468) <= dataBufferIn_long(2196);
	dataBufferOut_long(4211) <= dataBufferIn_long(2197);
	dataBufferOut_long(4954) <= dataBufferIn_long(2198);
	dataBufferOut_long(5697) <= dataBufferIn_long(2199);
	dataBufferOut_long( 296) <= dataBufferIn_long(2200);
	dataBufferOut_long(1039) <= dataBufferIn_long(2201);
	dataBufferOut_long(1782) <= dataBufferIn_long(2202);
	dataBufferOut_long(2525) <= dataBufferIn_long(2203);
	dataBufferOut_long(3268) <= dataBufferIn_long(2204);
	dataBufferOut_long(4011) <= dataBufferIn_long(2205);
	dataBufferOut_long(4754) <= dataBufferIn_long(2206);
	dataBufferOut_long(5497) <= dataBufferIn_long(2207);
	dataBufferOut_long(  96) <= dataBufferIn_long(2208);
	dataBufferOut_long( 839) <= dataBufferIn_long(2209);
	dataBufferOut_long(1582) <= dataBufferIn_long(2210);
	dataBufferOut_long(2325) <= dataBufferIn_long(2211);
	dataBufferOut_long(3068) <= dataBufferIn_long(2212);
	dataBufferOut_long(3811) <= dataBufferIn_long(2213);
	dataBufferOut_long(4554) <= dataBufferIn_long(2214);
	dataBufferOut_long(5297) <= dataBufferIn_long(2215);
	dataBufferOut_long(6040) <= dataBufferIn_long(2216);
	dataBufferOut_long( 639) <= dataBufferIn_long(2217);
	dataBufferOut_long(1382) <= dataBufferIn_long(2218);
	dataBufferOut_long(2125) <= dataBufferIn_long(2219);
	dataBufferOut_long(2868) <= dataBufferIn_long(2220);
	dataBufferOut_long(3611) <= dataBufferIn_long(2221);
	dataBufferOut_long(4354) <= dataBufferIn_long(2222);
	dataBufferOut_long(5097) <= dataBufferIn_long(2223);
	dataBufferOut_long(5840) <= dataBufferIn_long(2224);
	dataBufferOut_long( 439) <= dataBufferIn_long(2225);
	dataBufferOut_long(1182) <= dataBufferIn_long(2226);
	dataBufferOut_long(1925) <= dataBufferIn_long(2227);
	dataBufferOut_long(2668) <= dataBufferIn_long(2228);
	dataBufferOut_long(3411) <= dataBufferIn_long(2229);
	dataBufferOut_long(4154) <= dataBufferIn_long(2230);
	dataBufferOut_long(4897) <= dataBufferIn_long(2231);
	dataBufferOut_long(5640) <= dataBufferIn_long(2232);
	dataBufferOut_long( 239) <= dataBufferIn_long(2233);
	dataBufferOut_long( 982) <= dataBufferIn_long(2234);
	dataBufferOut_long(1725) <= dataBufferIn_long(2235);
	dataBufferOut_long(2468) <= dataBufferIn_long(2236);
	dataBufferOut_long(3211) <= dataBufferIn_long(2237);
	dataBufferOut_long(3954) <= dataBufferIn_long(2238);
	dataBufferOut_long(4697) <= dataBufferIn_long(2239);
	dataBufferOut_long(5440) <= dataBufferIn_long(2240);
	dataBufferOut_long(  39) <= dataBufferIn_long(2241);
	dataBufferOut_long( 782) <= dataBufferIn_long(2242);
	dataBufferOut_long(1525) <= dataBufferIn_long(2243);
	dataBufferOut_long(2268) <= dataBufferIn_long(2244);
	dataBufferOut_long(3011) <= dataBufferIn_long(2245);
	dataBufferOut_long(3754) <= dataBufferIn_long(2246);
	dataBufferOut_long(4497) <= dataBufferIn_long(2247);
	dataBufferOut_long(5240) <= dataBufferIn_long(2248);
	dataBufferOut_long(5983) <= dataBufferIn_long(2249);
	dataBufferOut_long( 582) <= dataBufferIn_long(2250);
	dataBufferOut_long(1325) <= dataBufferIn_long(2251);
	dataBufferOut_long(2068) <= dataBufferIn_long(2252);
	dataBufferOut_long(2811) <= dataBufferIn_long(2253);
	dataBufferOut_long(3554) <= dataBufferIn_long(2254);
	dataBufferOut_long(4297) <= dataBufferIn_long(2255);
	dataBufferOut_long(5040) <= dataBufferIn_long(2256);
	dataBufferOut_long(5783) <= dataBufferIn_long(2257);
	dataBufferOut_long( 382) <= dataBufferIn_long(2258);
	dataBufferOut_long(1125) <= dataBufferIn_long(2259);
	dataBufferOut_long(1868) <= dataBufferIn_long(2260);
	dataBufferOut_long(2611) <= dataBufferIn_long(2261);
	dataBufferOut_long(3354) <= dataBufferIn_long(2262);
	dataBufferOut_long(4097) <= dataBufferIn_long(2263);
	dataBufferOut_long(4840) <= dataBufferIn_long(2264);
	dataBufferOut_long(5583) <= dataBufferIn_long(2265);
	dataBufferOut_long( 182) <= dataBufferIn_long(2266);
	dataBufferOut_long( 925) <= dataBufferIn_long(2267);
	dataBufferOut_long(1668) <= dataBufferIn_long(2268);
	dataBufferOut_long(2411) <= dataBufferIn_long(2269);
	dataBufferOut_long(3154) <= dataBufferIn_long(2270);
	dataBufferOut_long(3897) <= dataBufferIn_long(2271);
	dataBufferOut_long(4640) <= dataBufferIn_long(2272);
	dataBufferOut_long(5383) <= dataBufferIn_long(2273);
	dataBufferOut_long(6126) <= dataBufferIn_long(2274);
	dataBufferOut_long( 725) <= dataBufferIn_long(2275);
	dataBufferOut_long(1468) <= dataBufferIn_long(2276);
	dataBufferOut_long(2211) <= dataBufferIn_long(2277);
	dataBufferOut_long(2954) <= dataBufferIn_long(2278);
	dataBufferOut_long(3697) <= dataBufferIn_long(2279);
	dataBufferOut_long(4440) <= dataBufferIn_long(2280);
	dataBufferOut_long(5183) <= dataBufferIn_long(2281);
	dataBufferOut_long(5926) <= dataBufferIn_long(2282);
	dataBufferOut_long( 525) <= dataBufferIn_long(2283);
	dataBufferOut_long(1268) <= dataBufferIn_long(2284);
	dataBufferOut_long(2011) <= dataBufferIn_long(2285);
	dataBufferOut_long(2754) <= dataBufferIn_long(2286);
	dataBufferOut_long(3497) <= dataBufferIn_long(2287);
	dataBufferOut_long(4240) <= dataBufferIn_long(2288);
	dataBufferOut_long(4983) <= dataBufferIn_long(2289);
	dataBufferOut_long(5726) <= dataBufferIn_long(2290);
	dataBufferOut_long( 325) <= dataBufferIn_long(2291);
	dataBufferOut_long(1068) <= dataBufferIn_long(2292);
	dataBufferOut_long(1811) <= dataBufferIn_long(2293);
	dataBufferOut_long(2554) <= dataBufferIn_long(2294);
	dataBufferOut_long(3297) <= dataBufferIn_long(2295);
	dataBufferOut_long(4040) <= dataBufferIn_long(2296);
	dataBufferOut_long(4783) <= dataBufferIn_long(2297);
	dataBufferOut_long(5526) <= dataBufferIn_long(2298);
	dataBufferOut_long( 125) <= dataBufferIn_long(2299);
	dataBufferOut_long( 868) <= dataBufferIn_long(2300);
	dataBufferOut_long(1611) <= dataBufferIn_long(2301);
	dataBufferOut_long(2354) <= dataBufferIn_long(2302);
	dataBufferOut_long(3097) <= dataBufferIn_long(2303);
	dataBufferOut_long(3840) <= dataBufferIn_long(2304);
	dataBufferOut_long(4583) <= dataBufferIn_long(2305);
	dataBufferOut_long(5326) <= dataBufferIn_long(2306);
	dataBufferOut_long(6069) <= dataBufferIn_long(2307);
	dataBufferOut_long( 668) <= dataBufferIn_long(2308);
	dataBufferOut_long(1411) <= dataBufferIn_long(2309);
	dataBufferOut_long(2154) <= dataBufferIn_long(2310);
	dataBufferOut_long(2897) <= dataBufferIn_long(2311);
	dataBufferOut_long(3640) <= dataBufferIn_long(2312);
	dataBufferOut_long(4383) <= dataBufferIn_long(2313);
	dataBufferOut_long(5126) <= dataBufferIn_long(2314);
	dataBufferOut_long(5869) <= dataBufferIn_long(2315);
	dataBufferOut_long( 468) <= dataBufferIn_long(2316);
	dataBufferOut_long(1211) <= dataBufferIn_long(2317);
	dataBufferOut_long(1954) <= dataBufferIn_long(2318);
	dataBufferOut_long(2697) <= dataBufferIn_long(2319);
	dataBufferOut_long(3440) <= dataBufferIn_long(2320);
	dataBufferOut_long(4183) <= dataBufferIn_long(2321);
	dataBufferOut_long(4926) <= dataBufferIn_long(2322);
	dataBufferOut_long(5669) <= dataBufferIn_long(2323);
	dataBufferOut_long( 268) <= dataBufferIn_long(2324);
	dataBufferOut_long(1011) <= dataBufferIn_long(2325);
	dataBufferOut_long(1754) <= dataBufferIn_long(2326);
	dataBufferOut_long(2497) <= dataBufferIn_long(2327);
	dataBufferOut_long(3240) <= dataBufferIn_long(2328);
	dataBufferOut_long(3983) <= dataBufferIn_long(2329);
	dataBufferOut_long(4726) <= dataBufferIn_long(2330);
	dataBufferOut_long(5469) <= dataBufferIn_long(2331);
	dataBufferOut_long(  68) <= dataBufferIn_long(2332);
	dataBufferOut_long( 811) <= dataBufferIn_long(2333);
	dataBufferOut_long(1554) <= dataBufferIn_long(2334);
	dataBufferOut_long(2297) <= dataBufferIn_long(2335);
	dataBufferOut_long(3040) <= dataBufferIn_long(2336);
	dataBufferOut_long(3783) <= dataBufferIn_long(2337);
	dataBufferOut_long(4526) <= dataBufferIn_long(2338);
	dataBufferOut_long(5269) <= dataBufferIn_long(2339);
	dataBufferOut_long(6012) <= dataBufferIn_long(2340);
	dataBufferOut_long( 611) <= dataBufferIn_long(2341);
	dataBufferOut_long(1354) <= dataBufferIn_long(2342);
	dataBufferOut_long(2097) <= dataBufferIn_long(2343);
	dataBufferOut_long(2840) <= dataBufferIn_long(2344);
	dataBufferOut_long(3583) <= dataBufferIn_long(2345);
	dataBufferOut_long(4326) <= dataBufferIn_long(2346);
	dataBufferOut_long(5069) <= dataBufferIn_long(2347);
	dataBufferOut_long(5812) <= dataBufferIn_long(2348);
	dataBufferOut_long( 411) <= dataBufferIn_long(2349);
	dataBufferOut_long(1154) <= dataBufferIn_long(2350);
	dataBufferOut_long(1897) <= dataBufferIn_long(2351);
	dataBufferOut_long(2640) <= dataBufferIn_long(2352);
	dataBufferOut_long(3383) <= dataBufferIn_long(2353);
	dataBufferOut_long(4126) <= dataBufferIn_long(2354);
	dataBufferOut_long(4869) <= dataBufferIn_long(2355);
	dataBufferOut_long(5612) <= dataBufferIn_long(2356);
	dataBufferOut_long( 211) <= dataBufferIn_long(2357);
	dataBufferOut_long( 954) <= dataBufferIn_long(2358);
	dataBufferOut_long(1697) <= dataBufferIn_long(2359);
	dataBufferOut_long(2440) <= dataBufferIn_long(2360);
	dataBufferOut_long(3183) <= dataBufferIn_long(2361);
	dataBufferOut_long(3926) <= dataBufferIn_long(2362);
	dataBufferOut_long(4669) <= dataBufferIn_long(2363);
	dataBufferOut_long(5412) <= dataBufferIn_long(2364);
	dataBufferOut_long(  11) <= dataBufferIn_long(2365);
	dataBufferOut_long( 754) <= dataBufferIn_long(2366);
	dataBufferOut_long(1497) <= dataBufferIn_long(2367);
	dataBufferOut_long(2240) <= dataBufferIn_long(2368);
	dataBufferOut_long(2983) <= dataBufferIn_long(2369);
	dataBufferOut_long(3726) <= dataBufferIn_long(2370);
	dataBufferOut_long(4469) <= dataBufferIn_long(2371);
	dataBufferOut_long(5212) <= dataBufferIn_long(2372);
	dataBufferOut_long(5955) <= dataBufferIn_long(2373);
	dataBufferOut_long( 554) <= dataBufferIn_long(2374);
	dataBufferOut_long(1297) <= dataBufferIn_long(2375);
	dataBufferOut_long(2040) <= dataBufferIn_long(2376);
	dataBufferOut_long(2783) <= dataBufferIn_long(2377);
	dataBufferOut_long(3526) <= dataBufferIn_long(2378);
	dataBufferOut_long(4269) <= dataBufferIn_long(2379);
	dataBufferOut_long(5012) <= dataBufferIn_long(2380);
	dataBufferOut_long(5755) <= dataBufferIn_long(2381);
	dataBufferOut_long( 354) <= dataBufferIn_long(2382);
	dataBufferOut_long(1097) <= dataBufferIn_long(2383);
	dataBufferOut_long(1840) <= dataBufferIn_long(2384);
	dataBufferOut_long(2583) <= dataBufferIn_long(2385);
	dataBufferOut_long(3326) <= dataBufferIn_long(2386);
	dataBufferOut_long(4069) <= dataBufferIn_long(2387);
	dataBufferOut_long(4812) <= dataBufferIn_long(2388);
	dataBufferOut_long(5555) <= dataBufferIn_long(2389);
	dataBufferOut_long( 154) <= dataBufferIn_long(2390);
	dataBufferOut_long( 897) <= dataBufferIn_long(2391);
	dataBufferOut_long(1640) <= dataBufferIn_long(2392);
	dataBufferOut_long(2383) <= dataBufferIn_long(2393);
	dataBufferOut_long(3126) <= dataBufferIn_long(2394);
	dataBufferOut_long(3869) <= dataBufferIn_long(2395);
	dataBufferOut_long(4612) <= dataBufferIn_long(2396);
	dataBufferOut_long(5355) <= dataBufferIn_long(2397);
	dataBufferOut_long(6098) <= dataBufferIn_long(2398);
	dataBufferOut_long( 697) <= dataBufferIn_long(2399);
	dataBufferOut_long(1440) <= dataBufferIn_long(2400);
	dataBufferOut_long(2183) <= dataBufferIn_long(2401);
	dataBufferOut_long(2926) <= dataBufferIn_long(2402);
	dataBufferOut_long(3669) <= dataBufferIn_long(2403);
	dataBufferOut_long(4412) <= dataBufferIn_long(2404);
	dataBufferOut_long(5155) <= dataBufferIn_long(2405);
	dataBufferOut_long(5898) <= dataBufferIn_long(2406);
	dataBufferOut_long( 497) <= dataBufferIn_long(2407);
	dataBufferOut_long(1240) <= dataBufferIn_long(2408);
	dataBufferOut_long(1983) <= dataBufferIn_long(2409);
	dataBufferOut_long(2726) <= dataBufferIn_long(2410);
	dataBufferOut_long(3469) <= dataBufferIn_long(2411);
	dataBufferOut_long(4212) <= dataBufferIn_long(2412);
	dataBufferOut_long(4955) <= dataBufferIn_long(2413);
	dataBufferOut_long(5698) <= dataBufferIn_long(2414);
	dataBufferOut_long( 297) <= dataBufferIn_long(2415);
	dataBufferOut_long(1040) <= dataBufferIn_long(2416);
	dataBufferOut_long(1783) <= dataBufferIn_long(2417);
	dataBufferOut_long(2526) <= dataBufferIn_long(2418);
	dataBufferOut_long(3269) <= dataBufferIn_long(2419);
	dataBufferOut_long(4012) <= dataBufferIn_long(2420);
	dataBufferOut_long(4755) <= dataBufferIn_long(2421);
	dataBufferOut_long(5498) <= dataBufferIn_long(2422);
	dataBufferOut_long(  97) <= dataBufferIn_long(2423);
	dataBufferOut_long( 840) <= dataBufferIn_long(2424);
	dataBufferOut_long(1583) <= dataBufferIn_long(2425);
	dataBufferOut_long(2326) <= dataBufferIn_long(2426);
	dataBufferOut_long(3069) <= dataBufferIn_long(2427);
	dataBufferOut_long(3812) <= dataBufferIn_long(2428);
	dataBufferOut_long(4555) <= dataBufferIn_long(2429);
	dataBufferOut_long(5298) <= dataBufferIn_long(2430);
	dataBufferOut_long(6041) <= dataBufferIn_long(2431);
	dataBufferOut_long( 640) <= dataBufferIn_long(2432);
	dataBufferOut_long(1383) <= dataBufferIn_long(2433);
	dataBufferOut_long(2126) <= dataBufferIn_long(2434);
	dataBufferOut_long(2869) <= dataBufferIn_long(2435);
	dataBufferOut_long(3612) <= dataBufferIn_long(2436);
	dataBufferOut_long(4355) <= dataBufferIn_long(2437);
	dataBufferOut_long(5098) <= dataBufferIn_long(2438);
	dataBufferOut_long(5841) <= dataBufferIn_long(2439);
	dataBufferOut_long( 440) <= dataBufferIn_long(2440);
	dataBufferOut_long(1183) <= dataBufferIn_long(2441);
	dataBufferOut_long(1926) <= dataBufferIn_long(2442);
	dataBufferOut_long(2669) <= dataBufferIn_long(2443);
	dataBufferOut_long(3412) <= dataBufferIn_long(2444);
	dataBufferOut_long(4155) <= dataBufferIn_long(2445);
	dataBufferOut_long(4898) <= dataBufferIn_long(2446);
	dataBufferOut_long(5641) <= dataBufferIn_long(2447);
	dataBufferOut_long( 240) <= dataBufferIn_long(2448);
	dataBufferOut_long( 983) <= dataBufferIn_long(2449);
	dataBufferOut_long(1726) <= dataBufferIn_long(2450);
	dataBufferOut_long(2469) <= dataBufferIn_long(2451);
	dataBufferOut_long(3212) <= dataBufferIn_long(2452);
	dataBufferOut_long(3955) <= dataBufferIn_long(2453);
	dataBufferOut_long(4698) <= dataBufferIn_long(2454);
	dataBufferOut_long(5441) <= dataBufferIn_long(2455);
	dataBufferOut_long(  40) <= dataBufferIn_long(2456);
	dataBufferOut_long( 783) <= dataBufferIn_long(2457);
	dataBufferOut_long(1526) <= dataBufferIn_long(2458);
	dataBufferOut_long(2269) <= dataBufferIn_long(2459);
	dataBufferOut_long(3012) <= dataBufferIn_long(2460);
	dataBufferOut_long(3755) <= dataBufferIn_long(2461);
	dataBufferOut_long(4498) <= dataBufferIn_long(2462);
	dataBufferOut_long(5241) <= dataBufferIn_long(2463);
	dataBufferOut_long(5984) <= dataBufferIn_long(2464);
	dataBufferOut_long( 583) <= dataBufferIn_long(2465);
	dataBufferOut_long(1326) <= dataBufferIn_long(2466);
	dataBufferOut_long(2069) <= dataBufferIn_long(2467);
	dataBufferOut_long(2812) <= dataBufferIn_long(2468);
	dataBufferOut_long(3555) <= dataBufferIn_long(2469);
	dataBufferOut_long(4298) <= dataBufferIn_long(2470);
	dataBufferOut_long(5041) <= dataBufferIn_long(2471);
	dataBufferOut_long(5784) <= dataBufferIn_long(2472);
	dataBufferOut_long( 383) <= dataBufferIn_long(2473);
	dataBufferOut_long(1126) <= dataBufferIn_long(2474);
	dataBufferOut_long(1869) <= dataBufferIn_long(2475);
	dataBufferOut_long(2612) <= dataBufferIn_long(2476);
	dataBufferOut_long(3355) <= dataBufferIn_long(2477);
	dataBufferOut_long(4098) <= dataBufferIn_long(2478);
	dataBufferOut_long(4841) <= dataBufferIn_long(2479);
	dataBufferOut_long(5584) <= dataBufferIn_long(2480);
	dataBufferOut_long( 183) <= dataBufferIn_long(2481);
	dataBufferOut_long( 926) <= dataBufferIn_long(2482);
	dataBufferOut_long(1669) <= dataBufferIn_long(2483);
	dataBufferOut_long(2412) <= dataBufferIn_long(2484);
	dataBufferOut_long(3155) <= dataBufferIn_long(2485);
	dataBufferOut_long(3898) <= dataBufferIn_long(2486);
	dataBufferOut_long(4641) <= dataBufferIn_long(2487);
	dataBufferOut_long(5384) <= dataBufferIn_long(2488);
	dataBufferOut_long(6127) <= dataBufferIn_long(2489);
	dataBufferOut_long( 726) <= dataBufferIn_long(2490);
	dataBufferOut_long(1469) <= dataBufferIn_long(2491);
	dataBufferOut_long(2212) <= dataBufferIn_long(2492);
	dataBufferOut_long(2955) <= dataBufferIn_long(2493);
	dataBufferOut_long(3698) <= dataBufferIn_long(2494);
	dataBufferOut_long(4441) <= dataBufferIn_long(2495);
	dataBufferOut_long(5184) <= dataBufferIn_long(2496);
	dataBufferOut_long(5927) <= dataBufferIn_long(2497);
	dataBufferOut_long( 526) <= dataBufferIn_long(2498);
	dataBufferOut_long(1269) <= dataBufferIn_long(2499);
	dataBufferOut_long(2012) <= dataBufferIn_long(2500);
	dataBufferOut_long(2755) <= dataBufferIn_long(2501);
	dataBufferOut_long(3498) <= dataBufferIn_long(2502);
	dataBufferOut_long(4241) <= dataBufferIn_long(2503);
	dataBufferOut_long(4984) <= dataBufferIn_long(2504);
	dataBufferOut_long(5727) <= dataBufferIn_long(2505);
	dataBufferOut_long( 326) <= dataBufferIn_long(2506);
	dataBufferOut_long(1069) <= dataBufferIn_long(2507);
	dataBufferOut_long(1812) <= dataBufferIn_long(2508);
	dataBufferOut_long(2555) <= dataBufferIn_long(2509);
	dataBufferOut_long(3298) <= dataBufferIn_long(2510);
	dataBufferOut_long(4041) <= dataBufferIn_long(2511);
	dataBufferOut_long(4784) <= dataBufferIn_long(2512);
	dataBufferOut_long(5527) <= dataBufferIn_long(2513);
	dataBufferOut_long( 126) <= dataBufferIn_long(2514);
	dataBufferOut_long( 869) <= dataBufferIn_long(2515);
	dataBufferOut_long(1612) <= dataBufferIn_long(2516);
	dataBufferOut_long(2355) <= dataBufferIn_long(2517);
	dataBufferOut_long(3098) <= dataBufferIn_long(2518);
	dataBufferOut_long(3841) <= dataBufferIn_long(2519);
	dataBufferOut_long(4584) <= dataBufferIn_long(2520);
	dataBufferOut_long(5327) <= dataBufferIn_long(2521);
	dataBufferOut_long(6070) <= dataBufferIn_long(2522);
	dataBufferOut_long( 669) <= dataBufferIn_long(2523);
	dataBufferOut_long(1412) <= dataBufferIn_long(2524);
	dataBufferOut_long(2155) <= dataBufferIn_long(2525);
	dataBufferOut_long(2898) <= dataBufferIn_long(2526);
	dataBufferOut_long(3641) <= dataBufferIn_long(2527);
	dataBufferOut_long(4384) <= dataBufferIn_long(2528);
	dataBufferOut_long(5127) <= dataBufferIn_long(2529);
	dataBufferOut_long(5870) <= dataBufferIn_long(2530);
	dataBufferOut_long( 469) <= dataBufferIn_long(2531);
	dataBufferOut_long(1212) <= dataBufferIn_long(2532);
	dataBufferOut_long(1955) <= dataBufferIn_long(2533);
	dataBufferOut_long(2698) <= dataBufferIn_long(2534);
	dataBufferOut_long(3441) <= dataBufferIn_long(2535);
	dataBufferOut_long(4184) <= dataBufferIn_long(2536);
	dataBufferOut_long(4927) <= dataBufferIn_long(2537);
	dataBufferOut_long(5670) <= dataBufferIn_long(2538);
	dataBufferOut_long( 269) <= dataBufferIn_long(2539);
	dataBufferOut_long(1012) <= dataBufferIn_long(2540);
	dataBufferOut_long(1755) <= dataBufferIn_long(2541);
	dataBufferOut_long(2498) <= dataBufferIn_long(2542);
	dataBufferOut_long(3241) <= dataBufferIn_long(2543);
	dataBufferOut_long(3984) <= dataBufferIn_long(2544);
	dataBufferOut_long(4727) <= dataBufferIn_long(2545);
	dataBufferOut_long(5470) <= dataBufferIn_long(2546);
	dataBufferOut_long(  69) <= dataBufferIn_long(2547);
	dataBufferOut_long( 812) <= dataBufferIn_long(2548);
	dataBufferOut_long(1555) <= dataBufferIn_long(2549);
	dataBufferOut_long(2298) <= dataBufferIn_long(2550);
	dataBufferOut_long(3041) <= dataBufferIn_long(2551);
	dataBufferOut_long(3784) <= dataBufferIn_long(2552);
	dataBufferOut_long(4527) <= dataBufferIn_long(2553);
	dataBufferOut_long(5270) <= dataBufferIn_long(2554);
	dataBufferOut_long(6013) <= dataBufferIn_long(2555);
	dataBufferOut_long( 612) <= dataBufferIn_long(2556);
	dataBufferOut_long(1355) <= dataBufferIn_long(2557);
	dataBufferOut_long(2098) <= dataBufferIn_long(2558);
	dataBufferOut_long(2841) <= dataBufferIn_long(2559);
	dataBufferOut_long(3584) <= dataBufferIn_long(2560);
	dataBufferOut_long(4327) <= dataBufferIn_long(2561);
	dataBufferOut_long(5070) <= dataBufferIn_long(2562);
	dataBufferOut_long(5813) <= dataBufferIn_long(2563);
	dataBufferOut_long( 412) <= dataBufferIn_long(2564);
	dataBufferOut_long(1155) <= dataBufferIn_long(2565);
	dataBufferOut_long(1898) <= dataBufferIn_long(2566);
	dataBufferOut_long(2641) <= dataBufferIn_long(2567);
	dataBufferOut_long(3384) <= dataBufferIn_long(2568);
	dataBufferOut_long(4127) <= dataBufferIn_long(2569);
	dataBufferOut_long(4870) <= dataBufferIn_long(2570);
	dataBufferOut_long(5613) <= dataBufferIn_long(2571);
	dataBufferOut_long( 212) <= dataBufferIn_long(2572);
	dataBufferOut_long( 955) <= dataBufferIn_long(2573);
	dataBufferOut_long(1698) <= dataBufferIn_long(2574);
	dataBufferOut_long(2441) <= dataBufferIn_long(2575);
	dataBufferOut_long(3184) <= dataBufferIn_long(2576);
	dataBufferOut_long(3927) <= dataBufferIn_long(2577);
	dataBufferOut_long(4670) <= dataBufferIn_long(2578);
	dataBufferOut_long(5413) <= dataBufferIn_long(2579);
	dataBufferOut_long(  12) <= dataBufferIn_long(2580);
	dataBufferOut_long( 755) <= dataBufferIn_long(2581);
	dataBufferOut_long(1498) <= dataBufferIn_long(2582);
	dataBufferOut_long(2241) <= dataBufferIn_long(2583);
	dataBufferOut_long(2984) <= dataBufferIn_long(2584);
	dataBufferOut_long(3727) <= dataBufferIn_long(2585);
	dataBufferOut_long(4470) <= dataBufferIn_long(2586);
	dataBufferOut_long(5213) <= dataBufferIn_long(2587);
	dataBufferOut_long(5956) <= dataBufferIn_long(2588);
	dataBufferOut_long( 555) <= dataBufferIn_long(2589);
	dataBufferOut_long(1298) <= dataBufferIn_long(2590);
	dataBufferOut_long(2041) <= dataBufferIn_long(2591);
	dataBufferOut_long(2784) <= dataBufferIn_long(2592);
	dataBufferOut_long(3527) <= dataBufferIn_long(2593);
	dataBufferOut_long(4270) <= dataBufferIn_long(2594);
	dataBufferOut_long(5013) <= dataBufferIn_long(2595);
	dataBufferOut_long(5756) <= dataBufferIn_long(2596);
	dataBufferOut_long( 355) <= dataBufferIn_long(2597);
	dataBufferOut_long(1098) <= dataBufferIn_long(2598);
	dataBufferOut_long(1841) <= dataBufferIn_long(2599);
	dataBufferOut_long(2584) <= dataBufferIn_long(2600);
	dataBufferOut_long(3327) <= dataBufferIn_long(2601);
	dataBufferOut_long(4070) <= dataBufferIn_long(2602);
	dataBufferOut_long(4813) <= dataBufferIn_long(2603);
	dataBufferOut_long(5556) <= dataBufferIn_long(2604);
	dataBufferOut_long( 155) <= dataBufferIn_long(2605);
	dataBufferOut_long( 898) <= dataBufferIn_long(2606);
	dataBufferOut_long(1641) <= dataBufferIn_long(2607);
	dataBufferOut_long(2384) <= dataBufferIn_long(2608);
	dataBufferOut_long(3127) <= dataBufferIn_long(2609);
	dataBufferOut_long(3870) <= dataBufferIn_long(2610);
	dataBufferOut_long(4613) <= dataBufferIn_long(2611);
	dataBufferOut_long(5356) <= dataBufferIn_long(2612);
	dataBufferOut_long(6099) <= dataBufferIn_long(2613);
	dataBufferOut_long( 698) <= dataBufferIn_long(2614);
	dataBufferOut_long(1441) <= dataBufferIn_long(2615);
	dataBufferOut_long(2184) <= dataBufferIn_long(2616);
	dataBufferOut_long(2927) <= dataBufferIn_long(2617);
	dataBufferOut_long(3670) <= dataBufferIn_long(2618);
	dataBufferOut_long(4413) <= dataBufferIn_long(2619);
	dataBufferOut_long(5156) <= dataBufferIn_long(2620);
	dataBufferOut_long(5899) <= dataBufferIn_long(2621);
	dataBufferOut_long( 498) <= dataBufferIn_long(2622);
	dataBufferOut_long(1241) <= dataBufferIn_long(2623);
	dataBufferOut_long(1984) <= dataBufferIn_long(2624);
	dataBufferOut_long(2727) <= dataBufferIn_long(2625);
	dataBufferOut_long(3470) <= dataBufferIn_long(2626);
	dataBufferOut_long(4213) <= dataBufferIn_long(2627);
	dataBufferOut_long(4956) <= dataBufferIn_long(2628);
	dataBufferOut_long(5699) <= dataBufferIn_long(2629);
	dataBufferOut_long( 298) <= dataBufferIn_long(2630);
	dataBufferOut_long(1041) <= dataBufferIn_long(2631);
	dataBufferOut_long(1784) <= dataBufferIn_long(2632);
	dataBufferOut_long(2527) <= dataBufferIn_long(2633);
	dataBufferOut_long(3270) <= dataBufferIn_long(2634);
	dataBufferOut_long(4013) <= dataBufferIn_long(2635);
	dataBufferOut_long(4756) <= dataBufferIn_long(2636);
	dataBufferOut_long(5499) <= dataBufferIn_long(2637);
	dataBufferOut_long(  98) <= dataBufferIn_long(2638);
	dataBufferOut_long( 841) <= dataBufferIn_long(2639);
	dataBufferOut_long(1584) <= dataBufferIn_long(2640);
	dataBufferOut_long(2327) <= dataBufferIn_long(2641);
	dataBufferOut_long(3070) <= dataBufferIn_long(2642);
	dataBufferOut_long(3813) <= dataBufferIn_long(2643);
	dataBufferOut_long(4556) <= dataBufferIn_long(2644);
	dataBufferOut_long(5299) <= dataBufferIn_long(2645);
	dataBufferOut_long(6042) <= dataBufferIn_long(2646);
	dataBufferOut_long( 641) <= dataBufferIn_long(2647);
	dataBufferOut_long(1384) <= dataBufferIn_long(2648);
	dataBufferOut_long(2127) <= dataBufferIn_long(2649);
	dataBufferOut_long(2870) <= dataBufferIn_long(2650);
	dataBufferOut_long(3613) <= dataBufferIn_long(2651);
	dataBufferOut_long(4356) <= dataBufferIn_long(2652);
	dataBufferOut_long(5099) <= dataBufferIn_long(2653);
	dataBufferOut_long(5842) <= dataBufferIn_long(2654);
	dataBufferOut_long( 441) <= dataBufferIn_long(2655);
	dataBufferOut_long(1184) <= dataBufferIn_long(2656);
	dataBufferOut_long(1927) <= dataBufferIn_long(2657);
	dataBufferOut_long(2670) <= dataBufferIn_long(2658);
	dataBufferOut_long(3413) <= dataBufferIn_long(2659);
	dataBufferOut_long(4156) <= dataBufferIn_long(2660);
	dataBufferOut_long(4899) <= dataBufferIn_long(2661);
	dataBufferOut_long(5642) <= dataBufferIn_long(2662);
	dataBufferOut_long( 241) <= dataBufferIn_long(2663);
	dataBufferOut_long( 984) <= dataBufferIn_long(2664);
	dataBufferOut_long(1727) <= dataBufferIn_long(2665);
	dataBufferOut_long(2470) <= dataBufferIn_long(2666);
	dataBufferOut_long(3213) <= dataBufferIn_long(2667);
	dataBufferOut_long(3956) <= dataBufferIn_long(2668);
	dataBufferOut_long(4699) <= dataBufferIn_long(2669);
	dataBufferOut_long(5442) <= dataBufferIn_long(2670);
	dataBufferOut_long(  41) <= dataBufferIn_long(2671);
	dataBufferOut_long( 784) <= dataBufferIn_long(2672);
	dataBufferOut_long(1527) <= dataBufferIn_long(2673);
	dataBufferOut_long(2270) <= dataBufferIn_long(2674);
	dataBufferOut_long(3013) <= dataBufferIn_long(2675);
	dataBufferOut_long(3756) <= dataBufferIn_long(2676);
	dataBufferOut_long(4499) <= dataBufferIn_long(2677);
	dataBufferOut_long(5242) <= dataBufferIn_long(2678);
	dataBufferOut_long(5985) <= dataBufferIn_long(2679);
	dataBufferOut_long( 584) <= dataBufferIn_long(2680);
	dataBufferOut_long(1327) <= dataBufferIn_long(2681);
	dataBufferOut_long(2070) <= dataBufferIn_long(2682);
	dataBufferOut_long(2813) <= dataBufferIn_long(2683);
	dataBufferOut_long(3556) <= dataBufferIn_long(2684);
	dataBufferOut_long(4299) <= dataBufferIn_long(2685);
	dataBufferOut_long(5042) <= dataBufferIn_long(2686);
	dataBufferOut_long(5785) <= dataBufferIn_long(2687);
	dataBufferOut_long( 384) <= dataBufferIn_long(2688);
	dataBufferOut_long(1127) <= dataBufferIn_long(2689);
	dataBufferOut_long(1870) <= dataBufferIn_long(2690);
	dataBufferOut_long(2613) <= dataBufferIn_long(2691);
	dataBufferOut_long(3356) <= dataBufferIn_long(2692);
	dataBufferOut_long(4099) <= dataBufferIn_long(2693);
	dataBufferOut_long(4842) <= dataBufferIn_long(2694);
	dataBufferOut_long(5585) <= dataBufferIn_long(2695);
	dataBufferOut_long( 184) <= dataBufferIn_long(2696);
	dataBufferOut_long( 927) <= dataBufferIn_long(2697);
	dataBufferOut_long(1670) <= dataBufferIn_long(2698);
	dataBufferOut_long(2413) <= dataBufferIn_long(2699);
	dataBufferOut_long(3156) <= dataBufferIn_long(2700);
	dataBufferOut_long(3899) <= dataBufferIn_long(2701);
	dataBufferOut_long(4642) <= dataBufferIn_long(2702);
	dataBufferOut_long(5385) <= dataBufferIn_long(2703);
	dataBufferOut_long(6128) <= dataBufferIn_long(2704);
	dataBufferOut_long( 727) <= dataBufferIn_long(2705);
	dataBufferOut_long(1470) <= dataBufferIn_long(2706);
	dataBufferOut_long(2213) <= dataBufferIn_long(2707);
	dataBufferOut_long(2956) <= dataBufferIn_long(2708);
	dataBufferOut_long(3699) <= dataBufferIn_long(2709);
	dataBufferOut_long(4442) <= dataBufferIn_long(2710);
	dataBufferOut_long(5185) <= dataBufferIn_long(2711);
	dataBufferOut_long(5928) <= dataBufferIn_long(2712);
	dataBufferOut_long( 527) <= dataBufferIn_long(2713);
	dataBufferOut_long(1270) <= dataBufferIn_long(2714);
	dataBufferOut_long(2013) <= dataBufferIn_long(2715);
	dataBufferOut_long(2756) <= dataBufferIn_long(2716);
	dataBufferOut_long(3499) <= dataBufferIn_long(2717);
	dataBufferOut_long(4242) <= dataBufferIn_long(2718);
	dataBufferOut_long(4985) <= dataBufferIn_long(2719);
	dataBufferOut_long(5728) <= dataBufferIn_long(2720);
	dataBufferOut_long( 327) <= dataBufferIn_long(2721);
	dataBufferOut_long(1070) <= dataBufferIn_long(2722);
	dataBufferOut_long(1813) <= dataBufferIn_long(2723);
	dataBufferOut_long(2556) <= dataBufferIn_long(2724);
	dataBufferOut_long(3299) <= dataBufferIn_long(2725);
	dataBufferOut_long(4042) <= dataBufferIn_long(2726);
	dataBufferOut_long(4785) <= dataBufferIn_long(2727);
	dataBufferOut_long(5528) <= dataBufferIn_long(2728);
	dataBufferOut_long( 127) <= dataBufferIn_long(2729);
	dataBufferOut_long( 870) <= dataBufferIn_long(2730);
	dataBufferOut_long(1613) <= dataBufferIn_long(2731);
	dataBufferOut_long(2356) <= dataBufferIn_long(2732);
	dataBufferOut_long(3099) <= dataBufferIn_long(2733);
	dataBufferOut_long(3842) <= dataBufferIn_long(2734);
	dataBufferOut_long(4585) <= dataBufferIn_long(2735);
	dataBufferOut_long(5328) <= dataBufferIn_long(2736);
	dataBufferOut_long(6071) <= dataBufferIn_long(2737);
	dataBufferOut_long( 670) <= dataBufferIn_long(2738);
	dataBufferOut_long(1413) <= dataBufferIn_long(2739);
	dataBufferOut_long(2156) <= dataBufferIn_long(2740);
	dataBufferOut_long(2899) <= dataBufferIn_long(2741);
	dataBufferOut_long(3642) <= dataBufferIn_long(2742);
	dataBufferOut_long(4385) <= dataBufferIn_long(2743);
	dataBufferOut_long(5128) <= dataBufferIn_long(2744);
	dataBufferOut_long(5871) <= dataBufferIn_long(2745);
	dataBufferOut_long( 470) <= dataBufferIn_long(2746);
	dataBufferOut_long(1213) <= dataBufferIn_long(2747);
	dataBufferOut_long(1956) <= dataBufferIn_long(2748);
	dataBufferOut_long(2699) <= dataBufferIn_long(2749);
	dataBufferOut_long(3442) <= dataBufferIn_long(2750);
	dataBufferOut_long(4185) <= dataBufferIn_long(2751);
	dataBufferOut_long(4928) <= dataBufferIn_long(2752);
	dataBufferOut_long(5671) <= dataBufferIn_long(2753);
	dataBufferOut_long( 270) <= dataBufferIn_long(2754);
	dataBufferOut_long(1013) <= dataBufferIn_long(2755);
	dataBufferOut_long(1756) <= dataBufferIn_long(2756);
	dataBufferOut_long(2499) <= dataBufferIn_long(2757);
	dataBufferOut_long(3242) <= dataBufferIn_long(2758);
	dataBufferOut_long(3985) <= dataBufferIn_long(2759);
	dataBufferOut_long(4728) <= dataBufferIn_long(2760);
	dataBufferOut_long(5471) <= dataBufferIn_long(2761);
	dataBufferOut_long(  70) <= dataBufferIn_long(2762);
	dataBufferOut_long( 813) <= dataBufferIn_long(2763);
	dataBufferOut_long(1556) <= dataBufferIn_long(2764);
	dataBufferOut_long(2299) <= dataBufferIn_long(2765);
	dataBufferOut_long(3042) <= dataBufferIn_long(2766);
	dataBufferOut_long(3785) <= dataBufferIn_long(2767);
	dataBufferOut_long(4528) <= dataBufferIn_long(2768);
	dataBufferOut_long(5271) <= dataBufferIn_long(2769);
	dataBufferOut_long(6014) <= dataBufferIn_long(2770);
	dataBufferOut_long( 613) <= dataBufferIn_long(2771);
	dataBufferOut_long(1356) <= dataBufferIn_long(2772);
	dataBufferOut_long(2099) <= dataBufferIn_long(2773);
	dataBufferOut_long(2842) <= dataBufferIn_long(2774);
	dataBufferOut_long(3585) <= dataBufferIn_long(2775);
	dataBufferOut_long(4328) <= dataBufferIn_long(2776);
	dataBufferOut_long(5071) <= dataBufferIn_long(2777);
	dataBufferOut_long(5814) <= dataBufferIn_long(2778);
	dataBufferOut_long( 413) <= dataBufferIn_long(2779);
	dataBufferOut_long(1156) <= dataBufferIn_long(2780);
	dataBufferOut_long(1899) <= dataBufferIn_long(2781);
	dataBufferOut_long(2642) <= dataBufferIn_long(2782);
	dataBufferOut_long(3385) <= dataBufferIn_long(2783);
	dataBufferOut_long(4128) <= dataBufferIn_long(2784);
	dataBufferOut_long(4871) <= dataBufferIn_long(2785);
	dataBufferOut_long(5614) <= dataBufferIn_long(2786);
	dataBufferOut_long( 213) <= dataBufferIn_long(2787);
	dataBufferOut_long( 956) <= dataBufferIn_long(2788);
	dataBufferOut_long(1699) <= dataBufferIn_long(2789);
	dataBufferOut_long(2442) <= dataBufferIn_long(2790);
	dataBufferOut_long(3185) <= dataBufferIn_long(2791);
	dataBufferOut_long(3928) <= dataBufferIn_long(2792);
	dataBufferOut_long(4671) <= dataBufferIn_long(2793);
	dataBufferOut_long(5414) <= dataBufferIn_long(2794);
	dataBufferOut_long(  13) <= dataBufferIn_long(2795);
	dataBufferOut_long( 756) <= dataBufferIn_long(2796);
	dataBufferOut_long(1499) <= dataBufferIn_long(2797);
	dataBufferOut_long(2242) <= dataBufferIn_long(2798);
	dataBufferOut_long(2985) <= dataBufferIn_long(2799);
	dataBufferOut_long(3728) <= dataBufferIn_long(2800);
	dataBufferOut_long(4471) <= dataBufferIn_long(2801);
	dataBufferOut_long(5214) <= dataBufferIn_long(2802);
	dataBufferOut_long(5957) <= dataBufferIn_long(2803);
	dataBufferOut_long( 556) <= dataBufferIn_long(2804);
	dataBufferOut_long(1299) <= dataBufferIn_long(2805);
	dataBufferOut_long(2042) <= dataBufferIn_long(2806);
	dataBufferOut_long(2785) <= dataBufferIn_long(2807);
	dataBufferOut_long(3528) <= dataBufferIn_long(2808);
	dataBufferOut_long(4271) <= dataBufferIn_long(2809);
	dataBufferOut_long(5014) <= dataBufferIn_long(2810);
	dataBufferOut_long(5757) <= dataBufferIn_long(2811);
	dataBufferOut_long( 356) <= dataBufferIn_long(2812);
	dataBufferOut_long(1099) <= dataBufferIn_long(2813);
	dataBufferOut_long(1842) <= dataBufferIn_long(2814);
	dataBufferOut_long(2585) <= dataBufferIn_long(2815);
	dataBufferOut_long(3328) <= dataBufferIn_long(2816);
	dataBufferOut_long(4071) <= dataBufferIn_long(2817);
	dataBufferOut_long(4814) <= dataBufferIn_long(2818);
	dataBufferOut_long(5557) <= dataBufferIn_long(2819);
	dataBufferOut_long( 156) <= dataBufferIn_long(2820);
	dataBufferOut_long( 899) <= dataBufferIn_long(2821);
	dataBufferOut_long(1642) <= dataBufferIn_long(2822);
	dataBufferOut_long(2385) <= dataBufferIn_long(2823);
	dataBufferOut_long(3128) <= dataBufferIn_long(2824);
	dataBufferOut_long(3871) <= dataBufferIn_long(2825);
	dataBufferOut_long(4614) <= dataBufferIn_long(2826);
	dataBufferOut_long(5357) <= dataBufferIn_long(2827);
	dataBufferOut_long(6100) <= dataBufferIn_long(2828);
	dataBufferOut_long( 699) <= dataBufferIn_long(2829);
	dataBufferOut_long(1442) <= dataBufferIn_long(2830);
	dataBufferOut_long(2185) <= dataBufferIn_long(2831);
	dataBufferOut_long(2928) <= dataBufferIn_long(2832);
	dataBufferOut_long(3671) <= dataBufferIn_long(2833);
	dataBufferOut_long(4414) <= dataBufferIn_long(2834);
	dataBufferOut_long(5157) <= dataBufferIn_long(2835);
	dataBufferOut_long(5900) <= dataBufferIn_long(2836);
	dataBufferOut_long( 499) <= dataBufferIn_long(2837);
	dataBufferOut_long(1242) <= dataBufferIn_long(2838);
	dataBufferOut_long(1985) <= dataBufferIn_long(2839);
	dataBufferOut_long(2728) <= dataBufferIn_long(2840);
	dataBufferOut_long(3471) <= dataBufferIn_long(2841);
	dataBufferOut_long(4214) <= dataBufferIn_long(2842);
	dataBufferOut_long(4957) <= dataBufferIn_long(2843);
	dataBufferOut_long(5700) <= dataBufferIn_long(2844);
	dataBufferOut_long( 299) <= dataBufferIn_long(2845);
	dataBufferOut_long(1042) <= dataBufferIn_long(2846);
	dataBufferOut_long(1785) <= dataBufferIn_long(2847);
	dataBufferOut_long(2528) <= dataBufferIn_long(2848);
	dataBufferOut_long(3271) <= dataBufferIn_long(2849);
	dataBufferOut_long(4014) <= dataBufferIn_long(2850);
	dataBufferOut_long(4757) <= dataBufferIn_long(2851);
	dataBufferOut_long(5500) <= dataBufferIn_long(2852);
	dataBufferOut_long(  99) <= dataBufferIn_long(2853);
	dataBufferOut_long( 842) <= dataBufferIn_long(2854);
	dataBufferOut_long(1585) <= dataBufferIn_long(2855);
	dataBufferOut_long(2328) <= dataBufferIn_long(2856);
	dataBufferOut_long(3071) <= dataBufferIn_long(2857);
	dataBufferOut_long(3814) <= dataBufferIn_long(2858);
	dataBufferOut_long(4557) <= dataBufferIn_long(2859);
	dataBufferOut_long(5300) <= dataBufferIn_long(2860);
	dataBufferOut_long(6043) <= dataBufferIn_long(2861);
	dataBufferOut_long( 642) <= dataBufferIn_long(2862);
	dataBufferOut_long(1385) <= dataBufferIn_long(2863);
	dataBufferOut_long(2128) <= dataBufferIn_long(2864);
	dataBufferOut_long(2871) <= dataBufferIn_long(2865);
	dataBufferOut_long(3614) <= dataBufferIn_long(2866);
	dataBufferOut_long(4357) <= dataBufferIn_long(2867);
	dataBufferOut_long(5100) <= dataBufferIn_long(2868);
	dataBufferOut_long(5843) <= dataBufferIn_long(2869);
	dataBufferOut_long( 442) <= dataBufferIn_long(2870);
	dataBufferOut_long(1185) <= dataBufferIn_long(2871);
	dataBufferOut_long(1928) <= dataBufferIn_long(2872);
	dataBufferOut_long(2671) <= dataBufferIn_long(2873);
	dataBufferOut_long(3414) <= dataBufferIn_long(2874);
	dataBufferOut_long(4157) <= dataBufferIn_long(2875);
	dataBufferOut_long(4900) <= dataBufferIn_long(2876);
	dataBufferOut_long(5643) <= dataBufferIn_long(2877);
	dataBufferOut_long( 242) <= dataBufferIn_long(2878);
	dataBufferOut_long( 985) <= dataBufferIn_long(2879);
	dataBufferOut_long(1728) <= dataBufferIn_long(2880);
	dataBufferOut_long(2471) <= dataBufferIn_long(2881);
	dataBufferOut_long(3214) <= dataBufferIn_long(2882);
	dataBufferOut_long(3957) <= dataBufferIn_long(2883);
	dataBufferOut_long(4700) <= dataBufferIn_long(2884);
	dataBufferOut_long(5443) <= dataBufferIn_long(2885);
	dataBufferOut_long(  42) <= dataBufferIn_long(2886);
	dataBufferOut_long( 785) <= dataBufferIn_long(2887);
	dataBufferOut_long(1528) <= dataBufferIn_long(2888);
	dataBufferOut_long(2271) <= dataBufferIn_long(2889);
	dataBufferOut_long(3014) <= dataBufferIn_long(2890);
	dataBufferOut_long(3757) <= dataBufferIn_long(2891);
	dataBufferOut_long(4500) <= dataBufferIn_long(2892);
	dataBufferOut_long(5243) <= dataBufferIn_long(2893);
	dataBufferOut_long(5986) <= dataBufferIn_long(2894);
	dataBufferOut_long( 585) <= dataBufferIn_long(2895);
	dataBufferOut_long(1328) <= dataBufferIn_long(2896);
	dataBufferOut_long(2071) <= dataBufferIn_long(2897);
	dataBufferOut_long(2814) <= dataBufferIn_long(2898);
	dataBufferOut_long(3557) <= dataBufferIn_long(2899);
	dataBufferOut_long(4300) <= dataBufferIn_long(2900);
	dataBufferOut_long(5043) <= dataBufferIn_long(2901);
	dataBufferOut_long(5786) <= dataBufferIn_long(2902);
	dataBufferOut_long( 385) <= dataBufferIn_long(2903);
	dataBufferOut_long(1128) <= dataBufferIn_long(2904);
	dataBufferOut_long(1871) <= dataBufferIn_long(2905);
	dataBufferOut_long(2614) <= dataBufferIn_long(2906);
	dataBufferOut_long(3357) <= dataBufferIn_long(2907);
	dataBufferOut_long(4100) <= dataBufferIn_long(2908);
	dataBufferOut_long(4843) <= dataBufferIn_long(2909);
	dataBufferOut_long(5586) <= dataBufferIn_long(2910);
	dataBufferOut_long( 185) <= dataBufferIn_long(2911);
	dataBufferOut_long( 928) <= dataBufferIn_long(2912);
	dataBufferOut_long(1671) <= dataBufferIn_long(2913);
	dataBufferOut_long(2414) <= dataBufferIn_long(2914);
	dataBufferOut_long(3157) <= dataBufferIn_long(2915);
	dataBufferOut_long(3900) <= dataBufferIn_long(2916);
	dataBufferOut_long(4643) <= dataBufferIn_long(2917);
	dataBufferOut_long(5386) <= dataBufferIn_long(2918);
	dataBufferOut_long(6129) <= dataBufferIn_long(2919);
	dataBufferOut_long( 728) <= dataBufferIn_long(2920);
	dataBufferOut_long(1471) <= dataBufferIn_long(2921);
	dataBufferOut_long(2214) <= dataBufferIn_long(2922);
	dataBufferOut_long(2957) <= dataBufferIn_long(2923);
	dataBufferOut_long(3700) <= dataBufferIn_long(2924);
	dataBufferOut_long(4443) <= dataBufferIn_long(2925);
	dataBufferOut_long(5186) <= dataBufferIn_long(2926);
	dataBufferOut_long(5929) <= dataBufferIn_long(2927);
	dataBufferOut_long( 528) <= dataBufferIn_long(2928);
	dataBufferOut_long(1271) <= dataBufferIn_long(2929);
	dataBufferOut_long(2014) <= dataBufferIn_long(2930);
	dataBufferOut_long(2757) <= dataBufferIn_long(2931);
	dataBufferOut_long(3500) <= dataBufferIn_long(2932);
	dataBufferOut_long(4243) <= dataBufferIn_long(2933);
	dataBufferOut_long(4986) <= dataBufferIn_long(2934);
	dataBufferOut_long(5729) <= dataBufferIn_long(2935);
	dataBufferOut_long( 328) <= dataBufferIn_long(2936);
	dataBufferOut_long(1071) <= dataBufferIn_long(2937);
	dataBufferOut_long(1814) <= dataBufferIn_long(2938);
	dataBufferOut_long(2557) <= dataBufferIn_long(2939);
	dataBufferOut_long(3300) <= dataBufferIn_long(2940);
	dataBufferOut_long(4043) <= dataBufferIn_long(2941);
	dataBufferOut_long(4786) <= dataBufferIn_long(2942);
	dataBufferOut_long(5529) <= dataBufferIn_long(2943);
	dataBufferOut_long( 128) <= dataBufferIn_long(2944);
	dataBufferOut_long( 871) <= dataBufferIn_long(2945);
	dataBufferOut_long(1614) <= dataBufferIn_long(2946);
	dataBufferOut_long(2357) <= dataBufferIn_long(2947);
	dataBufferOut_long(3100) <= dataBufferIn_long(2948);
	dataBufferOut_long(3843) <= dataBufferIn_long(2949);
	dataBufferOut_long(4586) <= dataBufferIn_long(2950);
	dataBufferOut_long(5329) <= dataBufferIn_long(2951);
	dataBufferOut_long(6072) <= dataBufferIn_long(2952);
	dataBufferOut_long( 671) <= dataBufferIn_long(2953);
	dataBufferOut_long(1414) <= dataBufferIn_long(2954);
	dataBufferOut_long(2157) <= dataBufferIn_long(2955);
	dataBufferOut_long(2900) <= dataBufferIn_long(2956);
	dataBufferOut_long(3643) <= dataBufferIn_long(2957);
	dataBufferOut_long(4386) <= dataBufferIn_long(2958);
	dataBufferOut_long(5129) <= dataBufferIn_long(2959);
	dataBufferOut_long(5872) <= dataBufferIn_long(2960);
	dataBufferOut_long( 471) <= dataBufferIn_long(2961);
	dataBufferOut_long(1214) <= dataBufferIn_long(2962);
	dataBufferOut_long(1957) <= dataBufferIn_long(2963);
	dataBufferOut_long(2700) <= dataBufferIn_long(2964);
	dataBufferOut_long(3443) <= dataBufferIn_long(2965);
	dataBufferOut_long(4186) <= dataBufferIn_long(2966);
	dataBufferOut_long(4929) <= dataBufferIn_long(2967);
	dataBufferOut_long(5672) <= dataBufferIn_long(2968);
	dataBufferOut_long( 271) <= dataBufferIn_long(2969);
	dataBufferOut_long(1014) <= dataBufferIn_long(2970);
	dataBufferOut_long(1757) <= dataBufferIn_long(2971);
	dataBufferOut_long(2500) <= dataBufferIn_long(2972);
	dataBufferOut_long(3243) <= dataBufferIn_long(2973);
	dataBufferOut_long(3986) <= dataBufferIn_long(2974);
	dataBufferOut_long(4729) <= dataBufferIn_long(2975);
	dataBufferOut_long(5472) <= dataBufferIn_long(2976);
	dataBufferOut_long(  71) <= dataBufferIn_long(2977);
	dataBufferOut_long( 814) <= dataBufferIn_long(2978);
	dataBufferOut_long(1557) <= dataBufferIn_long(2979);
	dataBufferOut_long(2300) <= dataBufferIn_long(2980);
	dataBufferOut_long(3043) <= dataBufferIn_long(2981);
	dataBufferOut_long(3786) <= dataBufferIn_long(2982);
	dataBufferOut_long(4529) <= dataBufferIn_long(2983);
	dataBufferOut_long(5272) <= dataBufferIn_long(2984);
	dataBufferOut_long(6015) <= dataBufferIn_long(2985);
	dataBufferOut_long( 614) <= dataBufferIn_long(2986);
	dataBufferOut_long(1357) <= dataBufferIn_long(2987);
	dataBufferOut_long(2100) <= dataBufferIn_long(2988);
	dataBufferOut_long(2843) <= dataBufferIn_long(2989);
	dataBufferOut_long(3586) <= dataBufferIn_long(2990);
	dataBufferOut_long(4329) <= dataBufferIn_long(2991);
	dataBufferOut_long(5072) <= dataBufferIn_long(2992);
	dataBufferOut_long(5815) <= dataBufferIn_long(2993);
	dataBufferOut_long( 414) <= dataBufferIn_long(2994);
	dataBufferOut_long(1157) <= dataBufferIn_long(2995);
	dataBufferOut_long(1900) <= dataBufferIn_long(2996);
	dataBufferOut_long(2643) <= dataBufferIn_long(2997);
	dataBufferOut_long(3386) <= dataBufferIn_long(2998);
	dataBufferOut_long(4129) <= dataBufferIn_long(2999);
	dataBufferOut_long(4872) <= dataBufferIn_long(3000);
	dataBufferOut_long(5615) <= dataBufferIn_long(3001);
	dataBufferOut_long( 214) <= dataBufferIn_long(3002);
	dataBufferOut_long( 957) <= dataBufferIn_long(3003);
	dataBufferOut_long(1700) <= dataBufferIn_long(3004);
	dataBufferOut_long(2443) <= dataBufferIn_long(3005);
	dataBufferOut_long(3186) <= dataBufferIn_long(3006);
	dataBufferOut_long(3929) <= dataBufferIn_long(3007);
	dataBufferOut_long(4672) <= dataBufferIn_long(3008);
	dataBufferOut_long(5415) <= dataBufferIn_long(3009);
	dataBufferOut_long(  14) <= dataBufferIn_long(3010);
	dataBufferOut_long( 757) <= dataBufferIn_long(3011);
	dataBufferOut_long(1500) <= dataBufferIn_long(3012);
	dataBufferOut_long(2243) <= dataBufferIn_long(3013);
	dataBufferOut_long(2986) <= dataBufferIn_long(3014);
	dataBufferOut_long(3729) <= dataBufferIn_long(3015);
	dataBufferOut_long(4472) <= dataBufferIn_long(3016);
	dataBufferOut_long(5215) <= dataBufferIn_long(3017);
	dataBufferOut_long(5958) <= dataBufferIn_long(3018);
	dataBufferOut_long( 557) <= dataBufferIn_long(3019);
	dataBufferOut_long(1300) <= dataBufferIn_long(3020);
	dataBufferOut_long(2043) <= dataBufferIn_long(3021);
	dataBufferOut_long(2786) <= dataBufferIn_long(3022);
	dataBufferOut_long(3529) <= dataBufferIn_long(3023);
	dataBufferOut_long(4272) <= dataBufferIn_long(3024);
	dataBufferOut_long(5015) <= dataBufferIn_long(3025);
	dataBufferOut_long(5758) <= dataBufferIn_long(3026);
	dataBufferOut_long( 357) <= dataBufferIn_long(3027);
	dataBufferOut_long(1100) <= dataBufferIn_long(3028);
	dataBufferOut_long(1843) <= dataBufferIn_long(3029);
	dataBufferOut_long(2586) <= dataBufferIn_long(3030);
	dataBufferOut_long(3329) <= dataBufferIn_long(3031);
	dataBufferOut_long(4072) <= dataBufferIn_long(3032);
	dataBufferOut_long(4815) <= dataBufferIn_long(3033);
	dataBufferOut_long(5558) <= dataBufferIn_long(3034);
	dataBufferOut_long( 157) <= dataBufferIn_long(3035);
	dataBufferOut_long( 900) <= dataBufferIn_long(3036);
	dataBufferOut_long(1643) <= dataBufferIn_long(3037);
	dataBufferOut_long(2386) <= dataBufferIn_long(3038);
	dataBufferOut_long(3129) <= dataBufferIn_long(3039);
	dataBufferOut_long(3872) <= dataBufferIn_long(3040);
	dataBufferOut_long(4615) <= dataBufferIn_long(3041);
	dataBufferOut_long(5358) <= dataBufferIn_long(3042);
	dataBufferOut_long(6101) <= dataBufferIn_long(3043);
	dataBufferOut_long( 700) <= dataBufferIn_long(3044);
	dataBufferOut_long(1443) <= dataBufferIn_long(3045);
	dataBufferOut_long(2186) <= dataBufferIn_long(3046);
	dataBufferOut_long(2929) <= dataBufferIn_long(3047);
	dataBufferOut_long(3672) <= dataBufferIn_long(3048);
	dataBufferOut_long(4415) <= dataBufferIn_long(3049);
	dataBufferOut_long(5158) <= dataBufferIn_long(3050);
	dataBufferOut_long(5901) <= dataBufferIn_long(3051);
	dataBufferOut_long( 500) <= dataBufferIn_long(3052);
	dataBufferOut_long(1243) <= dataBufferIn_long(3053);
	dataBufferOut_long(1986) <= dataBufferIn_long(3054);
	dataBufferOut_long(2729) <= dataBufferIn_long(3055);
	dataBufferOut_long(3472) <= dataBufferIn_long(3056);
	dataBufferOut_long(4215) <= dataBufferIn_long(3057);
	dataBufferOut_long(4958) <= dataBufferIn_long(3058);
	dataBufferOut_long(5701) <= dataBufferIn_long(3059);
	dataBufferOut_long( 300) <= dataBufferIn_long(3060);
	dataBufferOut_long(1043) <= dataBufferIn_long(3061);
	dataBufferOut_long(1786) <= dataBufferIn_long(3062);
	dataBufferOut_long(2529) <= dataBufferIn_long(3063);
	dataBufferOut_long(3272) <= dataBufferIn_long(3064);
	dataBufferOut_long(4015) <= dataBufferIn_long(3065);
	dataBufferOut_long(4758) <= dataBufferIn_long(3066);
	dataBufferOut_long(5501) <= dataBufferIn_long(3067);
	dataBufferOut_long( 100) <= dataBufferIn_long(3068);
	dataBufferOut_long( 843) <= dataBufferIn_long(3069);
	dataBufferOut_long(1586) <= dataBufferIn_long(3070);
	dataBufferOut_long(2329) <= dataBufferIn_long(3071);
	dataBufferOut_long(3072) <= dataBufferIn_long(3072);
	dataBufferOut_long(3815) <= dataBufferIn_long(3073);
	dataBufferOut_long(4558) <= dataBufferIn_long(3074);
	dataBufferOut_long(5301) <= dataBufferIn_long(3075);
	dataBufferOut_long(6044) <= dataBufferIn_long(3076);
	dataBufferOut_long( 643) <= dataBufferIn_long(3077);
	dataBufferOut_long(1386) <= dataBufferIn_long(3078);
	dataBufferOut_long(2129) <= dataBufferIn_long(3079);
	dataBufferOut_long(2872) <= dataBufferIn_long(3080);
	dataBufferOut_long(3615) <= dataBufferIn_long(3081);
	dataBufferOut_long(4358) <= dataBufferIn_long(3082);
	dataBufferOut_long(5101) <= dataBufferIn_long(3083);
	dataBufferOut_long(5844) <= dataBufferIn_long(3084);
	dataBufferOut_long( 443) <= dataBufferIn_long(3085);
	dataBufferOut_long(1186) <= dataBufferIn_long(3086);
	dataBufferOut_long(1929) <= dataBufferIn_long(3087);
	dataBufferOut_long(2672) <= dataBufferIn_long(3088);
	dataBufferOut_long(3415) <= dataBufferIn_long(3089);
	dataBufferOut_long(4158) <= dataBufferIn_long(3090);
	dataBufferOut_long(4901) <= dataBufferIn_long(3091);
	dataBufferOut_long(5644) <= dataBufferIn_long(3092);
	dataBufferOut_long( 243) <= dataBufferIn_long(3093);
	dataBufferOut_long( 986) <= dataBufferIn_long(3094);
	dataBufferOut_long(1729) <= dataBufferIn_long(3095);
	dataBufferOut_long(2472) <= dataBufferIn_long(3096);
	dataBufferOut_long(3215) <= dataBufferIn_long(3097);
	dataBufferOut_long(3958) <= dataBufferIn_long(3098);
	dataBufferOut_long(4701) <= dataBufferIn_long(3099);
	dataBufferOut_long(5444) <= dataBufferIn_long(3100);
	dataBufferOut_long(  43) <= dataBufferIn_long(3101);
	dataBufferOut_long( 786) <= dataBufferIn_long(3102);
	dataBufferOut_long(1529) <= dataBufferIn_long(3103);
	dataBufferOut_long(2272) <= dataBufferIn_long(3104);
	dataBufferOut_long(3015) <= dataBufferIn_long(3105);
	dataBufferOut_long(3758) <= dataBufferIn_long(3106);
	dataBufferOut_long(4501) <= dataBufferIn_long(3107);
	dataBufferOut_long(5244) <= dataBufferIn_long(3108);
	dataBufferOut_long(5987) <= dataBufferIn_long(3109);
	dataBufferOut_long( 586) <= dataBufferIn_long(3110);
	dataBufferOut_long(1329) <= dataBufferIn_long(3111);
	dataBufferOut_long(2072) <= dataBufferIn_long(3112);
	dataBufferOut_long(2815) <= dataBufferIn_long(3113);
	dataBufferOut_long(3558) <= dataBufferIn_long(3114);
	dataBufferOut_long(4301) <= dataBufferIn_long(3115);
	dataBufferOut_long(5044) <= dataBufferIn_long(3116);
	dataBufferOut_long(5787) <= dataBufferIn_long(3117);
	dataBufferOut_long( 386) <= dataBufferIn_long(3118);
	dataBufferOut_long(1129) <= dataBufferIn_long(3119);
	dataBufferOut_long(1872) <= dataBufferIn_long(3120);
	dataBufferOut_long(2615) <= dataBufferIn_long(3121);
	dataBufferOut_long(3358) <= dataBufferIn_long(3122);
	dataBufferOut_long(4101) <= dataBufferIn_long(3123);
	dataBufferOut_long(4844) <= dataBufferIn_long(3124);
	dataBufferOut_long(5587) <= dataBufferIn_long(3125);
	dataBufferOut_long( 186) <= dataBufferIn_long(3126);
	dataBufferOut_long( 929) <= dataBufferIn_long(3127);
	dataBufferOut_long(1672) <= dataBufferIn_long(3128);
	dataBufferOut_long(2415) <= dataBufferIn_long(3129);
	dataBufferOut_long(3158) <= dataBufferIn_long(3130);
	dataBufferOut_long(3901) <= dataBufferIn_long(3131);
	dataBufferOut_long(4644) <= dataBufferIn_long(3132);
	dataBufferOut_long(5387) <= dataBufferIn_long(3133);
	dataBufferOut_long(6130) <= dataBufferIn_long(3134);
	dataBufferOut_long( 729) <= dataBufferIn_long(3135);
	dataBufferOut_long(1472) <= dataBufferIn_long(3136);
	dataBufferOut_long(2215) <= dataBufferIn_long(3137);
	dataBufferOut_long(2958) <= dataBufferIn_long(3138);
	dataBufferOut_long(3701) <= dataBufferIn_long(3139);
	dataBufferOut_long(4444) <= dataBufferIn_long(3140);
	dataBufferOut_long(5187) <= dataBufferIn_long(3141);
	dataBufferOut_long(5930) <= dataBufferIn_long(3142);
	dataBufferOut_long( 529) <= dataBufferIn_long(3143);
	dataBufferOut_long(1272) <= dataBufferIn_long(3144);
	dataBufferOut_long(2015) <= dataBufferIn_long(3145);
	dataBufferOut_long(2758) <= dataBufferIn_long(3146);
	dataBufferOut_long(3501) <= dataBufferIn_long(3147);
	dataBufferOut_long(4244) <= dataBufferIn_long(3148);
	dataBufferOut_long(4987) <= dataBufferIn_long(3149);
	dataBufferOut_long(5730) <= dataBufferIn_long(3150);
	dataBufferOut_long( 329) <= dataBufferIn_long(3151);
	dataBufferOut_long(1072) <= dataBufferIn_long(3152);
	dataBufferOut_long(1815) <= dataBufferIn_long(3153);
	dataBufferOut_long(2558) <= dataBufferIn_long(3154);
	dataBufferOut_long(3301) <= dataBufferIn_long(3155);
	dataBufferOut_long(4044) <= dataBufferIn_long(3156);
	dataBufferOut_long(4787) <= dataBufferIn_long(3157);
	dataBufferOut_long(5530) <= dataBufferIn_long(3158);
	dataBufferOut_long( 129) <= dataBufferIn_long(3159);
	dataBufferOut_long( 872) <= dataBufferIn_long(3160);
	dataBufferOut_long(1615) <= dataBufferIn_long(3161);
	dataBufferOut_long(2358) <= dataBufferIn_long(3162);
	dataBufferOut_long(3101) <= dataBufferIn_long(3163);
	dataBufferOut_long(3844) <= dataBufferIn_long(3164);
	dataBufferOut_long(4587) <= dataBufferIn_long(3165);
	dataBufferOut_long(5330) <= dataBufferIn_long(3166);
	dataBufferOut_long(6073) <= dataBufferIn_long(3167);
	dataBufferOut_long( 672) <= dataBufferIn_long(3168);
	dataBufferOut_long(1415) <= dataBufferIn_long(3169);
	dataBufferOut_long(2158) <= dataBufferIn_long(3170);
	dataBufferOut_long(2901) <= dataBufferIn_long(3171);
	dataBufferOut_long(3644) <= dataBufferIn_long(3172);
	dataBufferOut_long(4387) <= dataBufferIn_long(3173);
	dataBufferOut_long(5130) <= dataBufferIn_long(3174);
	dataBufferOut_long(5873) <= dataBufferIn_long(3175);
	dataBufferOut_long( 472) <= dataBufferIn_long(3176);
	dataBufferOut_long(1215) <= dataBufferIn_long(3177);
	dataBufferOut_long(1958) <= dataBufferIn_long(3178);
	dataBufferOut_long(2701) <= dataBufferIn_long(3179);
	dataBufferOut_long(3444) <= dataBufferIn_long(3180);
	dataBufferOut_long(4187) <= dataBufferIn_long(3181);
	dataBufferOut_long(4930) <= dataBufferIn_long(3182);
	dataBufferOut_long(5673) <= dataBufferIn_long(3183);
	dataBufferOut_long( 272) <= dataBufferIn_long(3184);
	dataBufferOut_long(1015) <= dataBufferIn_long(3185);
	dataBufferOut_long(1758) <= dataBufferIn_long(3186);
	dataBufferOut_long(2501) <= dataBufferIn_long(3187);
	dataBufferOut_long(3244) <= dataBufferIn_long(3188);
	dataBufferOut_long(3987) <= dataBufferIn_long(3189);
	dataBufferOut_long(4730) <= dataBufferIn_long(3190);
	dataBufferOut_long(5473) <= dataBufferIn_long(3191);
	dataBufferOut_long(  72) <= dataBufferIn_long(3192);
	dataBufferOut_long( 815) <= dataBufferIn_long(3193);
	dataBufferOut_long(1558) <= dataBufferIn_long(3194);
	dataBufferOut_long(2301) <= dataBufferIn_long(3195);
	dataBufferOut_long(3044) <= dataBufferIn_long(3196);
	dataBufferOut_long(3787) <= dataBufferIn_long(3197);
	dataBufferOut_long(4530) <= dataBufferIn_long(3198);
	dataBufferOut_long(5273) <= dataBufferIn_long(3199);
	dataBufferOut_long(6016) <= dataBufferIn_long(3200);
	dataBufferOut_long( 615) <= dataBufferIn_long(3201);
	dataBufferOut_long(1358) <= dataBufferIn_long(3202);
	dataBufferOut_long(2101) <= dataBufferIn_long(3203);
	dataBufferOut_long(2844) <= dataBufferIn_long(3204);
	dataBufferOut_long(3587) <= dataBufferIn_long(3205);
	dataBufferOut_long(4330) <= dataBufferIn_long(3206);
	dataBufferOut_long(5073) <= dataBufferIn_long(3207);
	dataBufferOut_long(5816) <= dataBufferIn_long(3208);
	dataBufferOut_long( 415) <= dataBufferIn_long(3209);
	dataBufferOut_long(1158) <= dataBufferIn_long(3210);
	dataBufferOut_long(1901) <= dataBufferIn_long(3211);
	dataBufferOut_long(2644) <= dataBufferIn_long(3212);
	dataBufferOut_long(3387) <= dataBufferIn_long(3213);
	dataBufferOut_long(4130) <= dataBufferIn_long(3214);
	dataBufferOut_long(4873) <= dataBufferIn_long(3215);
	dataBufferOut_long(5616) <= dataBufferIn_long(3216);
	dataBufferOut_long( 215) <= dataBufferIn_long(3217);
	dataBufferOut_long( 958) <= dataBufferIn_long(3218);
	dataBufferOut_long(1701) <= dataBufferIn_long(3219);
	dataBufferOut_long(2444) <= dataBufferIn_long(3220);
	dataBufferOut_long(3187) <= dataBufferIn_long(3221);
	dataBufferOut_long(3930) <= dataBufferIn_long(3222);
	dataBufferOut_long(4673) <= dataBufferIn_long(3223);
	dataBufferOut_long(5416) <= dataBufferIn_long(3224);
	dataBufferOut_long(  15) <= dataBufferIn_long(3225);
	dataBufferOut_long( 758) <= dataBufferIn_long(3226);
	dataBufferOut_long(1501) <= dataBufferIn_long(3227);
	dataBufferOut_long(2244) <= dataBufferIn_long(3228);
	dataBufferOut_long(2987) <= dataBufferIn_long(3229);
	dataBufferOut_long(3730) <= dataBufferIn_long(3230);
	dataBufferOut_long(4473) <= dataBufferIn_long(3231);
	dataBufferOut_long(5216) <= dataBufferIn_long(3232);
	dataBufferOut_long(5959) <= dataBufferIn_long(3233);
	dataBufferOut_long( 558) <= dataBufferIn_long(3234);
	dataBufferOut_long(1301) <= dataBufferIn_long(3235);
	dataBufferOut_long(2044) <= dataBufferIn_long(3236);
	dataBufferOut_long(2787) <= dataBufferIn_long(3237);
	dataBufferOut_long(3530) <= dataBufferIn_long(3238);
	dataBufferOut_long(4273) <= dataBufferIn_long(3239);
	dataBufferOut_long(5016) <= dataBufferIn_long(3240);
	dataBufferOut_long(5759) <= dataBufferIn_long(3241);
	dataBufferOut_long( 358) <= dataBufferIn_long(3242);
	dataBufferOut_long(1101) <= dataBufferIn_long(3243);
	dataBufferOut_long(1844) <= dataBufferIn_long(3244);
	dataBufferOut_long(2587) <= dataBufferIn_long(3245);
	dataBufferOut_long(3330) <= dataBufferIn_long(3246);
	dataBufferOut_long(4073) <= dataBufferIn_long(3247);
	dataBufferOut_long(4816) <= dataBufferIn_long(3248);
	dataBufferOut_long(5559) <= dataBufferIn_long(3249);
	dataBufferOut_long( 158) <= dataBufferIn_long(3250);
	dataBufferOut_long( 901) <= dataBufferIn_long(3251);
	dataBufferOut_long(1644) <= dataBufferIn_long(3252);
	dataBufferOut_long(2387) <= dataBufferIn_long(3253);
	dataBufferOut_long(3130) <= dataBufferIn_long(3254);
	dataBufferOut_long(3873) <= dataBufferIn_long(3255);
	dataBufferOut_long(4616) <= dataBufferIn_long(3256);
	dataBufferOut_long(5359) <= dataBufferIn_long(3257);
	dataBufferOut_long(6102) <= dataBufferIn_long(3258);
	dataBufferOut_long( 701) <= dataBufferIn_long(3259);
	dataBufferOut_long(1444) <= dataBufferIn_long(3260);
	dataBufferOut_long(2187) <= dataBufferIn_long(3261);
	dataBufferOut_long(2930) <= dataBufferIn_long(3262);
	dataBufferOut_long(3673) <= dataBufferIn_long(3263);
	dataBufferOut_long(4416) <= dataBufferIn_long(3264);
	dataBufferOut_long(5159) <= dataBufferIn_long(3265);
	dataBufferOut_long(5902) <= dataBufferIn_long(3266);
	dataBufferOut_long( 501) <= dataBufferIn_long(3267);
	dataBufferOut_long(1244) <= dataBufferIn_long(3268);
	dataBufferOut_long(1987) <= dataBufferIn_long(3269);
	dataBufferOut_long(2730) <= dataBufferIn_long(3270);
	dataBufferOut_long(3473) <= dataBufferIn_long(3271);
	dataBufferOut_long(4216) <= dataBufferIn_long(3272);
	dataBufferOut_long(4959) <= dataBufferIn_long(3273);
	dataBufferOut_long(5702) <= dataBufferIn_long(3274);
	dataBufferOut_long( 301) <= dataBufferIn_long(3275);
	dataBufferOut_long(1044) <= dataBufferIn_long(3276);
	dataBufferOut_long(1787) <= dataBufferIn_long(3277);
	dataBufferOut_long(2530) <= dataBufferIn_long(3278);
	dataBufferOut_long(3273) <= dataBufferIn_long(3279);
	dataBufferOut_long(4016) <= dataBufferIn_long(3280);
	dataBufferOut_long(4759) <= dataBufferIn_long(3281);
	dataBufferOut_long(5502) <= dataBufferIn_long(3282);
	dataBufferOut_long( 101) <= dataBufferIn_long(3283);
	dataBufferOut_long( 844) <= dataBufferIn_long(3284);
	dataBufferOut_long(1587) <= dataBufferIn_long(3285);
	dataBufferOut_long(2330) <= dataBufferIn_long(3286);
	dataBufferOut_long(3073) <= dataBufferIn_long(3287);
	dataBufferOut_long(3816) <= dataBufferIn_long(3288);
	dataBufferOut_long(4559) <= dataBufferIn_long(3289);
	dataBufferOut_long(5302) <= dataBufferIn_long(3290);
	dataBufferOut_long(6045) <= dataBufferIn_long(3291);
	dataBufferOut_long( 644) <= dataBufferIn_long(3292);
	dataBufferOut_long(1387) <= dataBufferIn_long(3293);
	dataBufferOut_long(2130) <= dataBufferIn_long(3294);
	dataBufferOut_long(2873) <= dataBufferIn_long(3295);
	dataBufferOut_long(3616) <= dataBufferIn_long(3296);
	dataBufferOut_long(4359) <= dataBufferIn_long(3297);
	dataBufferOut_long(5102) <= dataBufferIn_long(3298);
	dataBufferOut_long(5845) <= dataBufferIn_long(3299);
	dataBufferOut_long( 444) <= dataBufferIn_long(3300);
	dataBufferOut_long(1187) <= dataBufferIn_long(3301);
	dataBufferOut_long(1930) <= dataBufferIn_long(3302);
	dataBufferOut_long(2673) <= dataBufferIn_long(3303);
	dataBufferOut_long(3416) <= dataBufferIn_long(3304);
	dataBufferOut_long(4159) <= dataBufferIn_long(3305);
	dataBufferOut_long(4902) <= dataBufferIn_long(3306);
	dataBufferOut_long(5645) <= dataBufferIn_long(3307);
	dataBufferOut_long( 244) <= dataBufferIn_long(3308);
	dataBufferOut_long( 987) <= dataBufferIn_long(3309);
	dataBufferOut_long(1730) <= dataBufferIn_long(3310);
	dataBufferOut_long(2473) <= dataBufferIn_long(3311);
	dataBufferOut_long(3216) <= dataBufferIn_long(3312);
	dataBufferOut_long(3959) <= dataBufferIn_long(3313);
	dataBufferOut_long(4702) <= dataBufferIn_long(3314);
	dataBufferOut_long(5445) <= dataBufferIn_long(3315);
	dataBufferOut_long(  44) <= dataBufferIn_long(3316);
	dataBufferOut_long( 787) <= dataBufferIn_long(3317);
	dataBufferOut_long(1530) <= dataBufferIn_long(3318);
	dataBufferOut_long(2273) <= dataBufferIn_long(3319);
	dataBufferOut_long(3016) <= dataBufferIn_long(3320);
	dataBufferOut_long(3759) <= dataBufferIn_long(3321);
	dataBufferOut_long(4502) <= dataBufferIn_long(3322);
	dataBufferOut_long(5245) <= dataBufferIn_long(3323);
	dataBufferOut_long(5988) <= dataBufferIn_long(3324);
	dataBufferOut_long( 587) <= dataBufferIn_long(3325);
	dataBufferOut_long(1330) <= dataBufferIn_long(3326);
	dataBufferOut_long(2073) <= dataBufferIn_long(3327);
	dataBufferOut_long(2816) <= dataBufferIn_long(3328);
	dataBufferOut_long(3559) <= dataBufferIn_long(3329);
	dataBufferOut_long(4302) <= dataBufferIn_long(3330);
	dataBufferOut_long(5045) <= dataBufferIn_long(3331);
	dataBufferOut_long(5788) <= dataBufferIn_long(3332);
	dataBufferOut_long( 387) <= dataBufferIn_long(3333);
	dataBufferOut_long(1130) <= dataBufferIn_long(3334);
	dataBufferOut_long(1873) <= dataBufferIn_long(3335);
	dataBufferOut_long(2616) <= dataBufferIn_long(3336);
	dataBufferOut_long(3359) <= dataBufferIn_long(3337);
	dataBufferOut_long(4102) <= dataBufferIn_long(3338);
	dataBufferOut_long(4845) <= dataBufferIn_long(3339);
	dataBufferOut_long(5588) <= dataBufferIn_long(3340);
	dataBufferOut_long( 187) <= dataBufferIn_long(3341);
	dataBufferOut_long( 930) <= dataBufferIn_long(3342);
	dataBufferOut_long(1673) <= dataBufferIn_long(3343);
	dataBufferOut_long(2416) <= dataBufferIn_long(3344);
	dataBufferOut_long(3159) <= dataBufferIn_long(3345);
	dataBufferOut_long(3902) <= dataBufferIn_long(3346);
	dataBufferOut_long(4645) <= dataBufferIn_long(3347);
	dataBufferOut_long(5388) <= dataBufferIn_long(3348);
	dataBufferOut_long(6131) <= dataBufferIn_long(3349);
	dataBufferOut_long( 730) <= dataBufferIn_long(3350);
	dataBufferOut_long(1473) <= dataBufferIn_long(3351);
	dataBufferOut_long(2216) <= dataBufferIn_long(3352);
	dataBufferOut_long(2959) <= dataBufferIn_long(3353);
	dataBufferOut_long(3702) <= dataBufferIn_long(3354);
	dataBufferOut_long(4445) <= dataBufferIn_long(3355);
	dataBufferOut_long(5188) <= dataBufferIn_long(3356);
	dataBufferOut_long(5931) <= dataBufferIn_long(3357);
	dataBufferOut_long( 530) <= dataBufferIn_long(3358);
	dataBufferOut_long(1273) <= dataBufferIn_long(3359);
	dataBufferOut_long(2016) <= dataBufferIn_long(3360);
	dataBufferOut_long(2759) <= dataBufferIn_long(3361);
	dataBufferOut_long(3502) <= dataBufferIn_long(3362);
	dataBufferOut_long(4245) <= dataBufferIn_long(3363);
	dataBufferOut_long(4988) <= dataBufferIn_long(3364);
	dataBufferOut_long(5731) <= dataBufferIn_long(3365);
	dataBufferOut_long( 330) <= dataBufferIn_long(3366);
	dataBufferOut_long(1073) <= dataBufferIn_long(3367);
	dataBufferOut_long(1816) <= dataBufferIn_long(3368);
	dataBufferOut_long(2559) <= dataBufferIn_long(3369);
	dataBufferOut_long(3302) <= dataBufferIn_long(3370);
	dataBufferOut_long(4045) <= dataBufferIn_long(3371);
	dataBufferOut_long(4788) <= dataBufferIn_long(3372);
	dataBufferOut_long(5531) <= dataBufferIn_long(3373);
	dataBufferOut_long( 130) <= dataBufferIn_long(3374);
	dataBufferOut_long( 873) <= dataBufferIn_long(3375);
	dataBufferOut_long(1616) <= dataBufferIn_long(3376);
	dataBufferOut_long(2359) <= dataBufferIn_long(3377);
	dataBufferOut_long(3102) <= dataBufferIn_long(3378);
	dataBufferOut_long(3845) <= dataBufferIn_long(3379);
	dataBufferOut_long(4588) <= dataBufferIn_long(3380);
	dataBufferOut_long(5331) <= dataBufferIn_long(3381);
	dataBufferOut_long(6074) <= dataBufferIn_long(3382);
	dataBufferOut_long( 673) <= dataBufferIn_long(3383);
	dataBufferOut_long(1416) <= dataBufferIn_long(3384);
	dataBufferOut_long(2159) <= dataBufferIn_long(3385);
	dataBufferOut_long(2902) <= dataBufferIn_long(3386);
	dataBufferOut_long(3645) <= dataBufferIn_long(3387);
	dataBufferOut_long(4388) <= dataBufferIn_long(3388);
	dataBufferOut_long(5131) <= dataBufferIn_long(3389);
	dataBufferOut_long(5874) <= dataBufferIn_long(3390);
	dataBufferOut_long( 473) <= dataBufferIn_long(3391);
	dataBufferOut_long(1216) <= dataBufferIn_long(3392);
	dataBufferOut_long(1959) <= dataBufferIn_long(3393);
	dataBufferOut_long(2702) <= dataBufferIn_long(3394);
	dataBufferOut_long(3445) <= dataBufferIn_long(3395);
	dataBufferOut_long(4188) <= dataBufferIn_long(3396);
	dataBufferOut_long(4931) <= dataBufferIn_long(3397);
	dataBufferOut_long(5674) <= dataBufferIn_long(3398);
	dataBufferOut_long( 273) <= dataBufferIn_long(3399);
	dataBufferOut_long(1016) <= dataBufferIn_long(3400);
	dataBufferOut_long(1759) <= dataBufferIn_long(3401);
	dataBufferOut_long(2502) <= dataBufferIn_long(3402);
	dataBufferOut_long(3245) <= dataBufferIn_long(3403);
	dataBufferOut_long(3988) <= dataBufferIn_long(3404);
	dataBufferOut_long(4731) <= dataBufferIn_long(3405);
	dataBufferOut_long(5474) <= dataBufferIn_long(3406);
	dataBufferOut_long(  73) <= dataBufferIn_long(3407);
	dataBufferOut_long( 816) <= dataBufferIn_long(3408);
	dataBufferOut_long(1559) <= dataBufferIn_long(3409);
	dataBufferOut_long(2302) <= dataBufferIn_long(3410);
	dataBufferOut_long(3045) <= dataBufferIn_long(3411);
	dataBufferOut_long(3788) <= dataBufferIn_long(3412);
	dataBufferOut_long(4531) <= dataBufferIn_long(3413);
	dataBufferOut_long(5274) <= dataBufferIn_long(3414);
	dataBufferOut_long(6017) <= dataBufferIn_long(3415);
	dataBufferOut_long( 616) <= dataBufferIn_long(3416);
	dataBufferOut_long(1359) <= dataBufferIn_long(3417);
	dataBufferOut_long(2102) <= dataBufferIn_long(3418);
	dataBufferOut_long(2845) <= dataBufferIn_long(3419);
	dataBufferOut_long(3588) <= dataBufferIn_long(3420);
	dataBufferOut_long(4331) <= dataBufferIn_long(3421);
	dataBufferOut_long(5074) <= dataBufferIn_long(3422);
	dataBufferOut_long(5817) <= dataBufferIn_long(3423);
	dataBufferOut_long( 416) <= dataBufferIn_long(3424);
	dataBufferOut_long(1159) <= dataBufferIn_long(3425);
	dataBufferOut_long(1902) <= dataBufferIn_long(3426);
	dataBufferOut_long(2645) <= dataBufferIn_long(3427);
	dataBufferOut_long(3388) <= dataBufferIn_long(3428);
	dataBufferOut_long(4131) <= dataBufferIn_long(3429);
	dataBufferOut_long(4874) <= dataBufferIn_long(3430);
	dataBufferOut_long(5617) <= dataBufferIn_long(3431);
	dataBufferOut_long( 216) <= dataBufferIn_long(3432);
	dataBufferOut_long( 959) <= dataBufferIn_long(3433);
	dataBufferOut_long(1702) <= dataBufferIn_long(3434);
	dataBufferOut_long(2445) <= dataBufferIn_long(3435);
	dataBufferOut_long(3188) <= dataBufferIn_long(3436);
	dataBufferOut_long(3931) <= dataBufferIn_long(3437);
	dataBufferOut_long(4674) <= dataBufferIn_long(3438);
	dataBufferOut_long(5417) <= dataBufferIn_long(3439);
	dataBufferOut_long(  16) <= dataBufferIn_long(3440);
	dataBufferOut_long( 759) <= dataBufferIn_long(3441);
	dataBufferOut_long(1502) <= dataBufferIn_long(3442);
	dataBufferOut_long(2245) <= dataBufferIn_long(3443);
	dataBufferOut_long(2988) <= dataBufferIn_long(3444);
	dataBufferOut_long(3731) <= dataBufferIn_long(3445);
	dataBufferOut_long(4474) <= dataBufferIn_long(3446);
	dataBufferOut_long(5217) <= dataBufferIn_long(3447);
	dataBufferOut_long(5960) <= dataBufferIn_long(3448);
	dataBufferOut_long( 559) <= dataBufferIn_long(3449);
	dataBufferOut_long(1302) <= dataBufferIn_long(3450);
	dataBufferOut_long(2045) <= dataBufferIn_long(3451);
	dataBufferOut_long(2788) <= dataBufferIn_long(3452);
	dataBufferOut_long(3531) <= dataBufferIn_long(3453);
	dataBufferOut_long(4274) <= dataBufferIn_long(3454);
	dataBufferOut_long(5017) <= dataBufferIn_long(3455);
	dataBufferOut_long(5760) <= dataBufferIn_long(3456);
	dataBufferOut_long( 359) <= dataBufferIn_long(3457);
	dataBufferOut_long(1102) <= dataBufferIn_long(3458);
	dataBufferOut_long(1845) <= dataBufferIn_long(3459);
	dataBufferOut_long(2588) <= dataBufferIn_long(3460);
	dataBufferOut_long(3331) <= dataBufferIn_long(3461);
	dataBufferOut_long(4074) <= dataBufferIn_long(3462);
	dataBufferOut_long(4817) <= dataBufferIn_long(3463);
	dataBufferOut_long(5560) <= dataBufferIn_long(3464);
	dataBufferOut_long( 159) <= dataBufferIn_long(3465);
	dataBufferOut_long( 902) <= dataBufferIn_long(3466);
	dataBufferOut_long(1645) <= dataBufferIn_long(3467);
	dataBufferOut_long(2388) <= dataBufferIn_long(3468);
	dataBufferOut_long(3131) <= dataBufferIn_long(3469);
	dataBufferOut_long(3874) <= dataBufferIn_long(3470);
	dataBufferOut_long(4617) <= dataBufferIn_long(3471);
	dataBufferOut_long(5360) <= dataBufferIn_long(3472);
	dataBufferOut_long(6103) <= dataBufferIn_long(3473);
	dataBufferOut_long( 702) <= dataBufferIn_long(3474);
	dataBufferOut_long(1445) <= dataBufferIn_long(3475);
	dataBufferOut_long(2188) <= dataBufferIn_long(3476);
	dataBufferOut_long(2931) <= dataBufferIn_long(3477);
	dataBufferOut_long(3674) <= dataBufferIn_long(3478);
	dataBufferOut_long(4417) <= dataBufferIn_long(3479);
	dataBufferOut_long(5160) <= dataBufferIn_long(3480);
	dataBufferOut_long(5903) <= dataBufferIn_long(3481);
	dataBufferOut_long( 502) <= dataBufferIn_long(3482);
	dataBufferOut_long(1245) <= dataBufferIn_long(3483);
	dataBufferOut_long(1988) <= dataBufferIn_long(3484);
	dataBufferOut_long(2731) <= dataBufferIn_long(3485);
	dataBufferOut_long(3474) <= dataBufferIn_long(3486);
	dataBufferOut_long(4217) <= dataBufferIn_long(3487);
	dataBufferOut_long(4960) <= dataBufferIn_long(3488);
	dataBufferOut_long(5703) <= dataBufferIn_long(3489);
	dataBufferOut_long( 302) <= dataBufferIn_long(3490);
	dataBufferOut_long(1045) <= dataBufferIn_long(3491);
	dataBufferOut_long(1788) <= dataBufferIn_long(3492);
	dataBufferOut_long(2531) <= dataBufferIn_long(3493);
	dataBufferOut_long(3274) <= dataBufferIn_long(3494);
	dataBufferOut_long(4017) <= dataBufferIn_long(3495);
	dataBufferOut_long(4760) <= dataBufferIn_long(3496);
	dataBufferOut_long(5503) <= dataBufferIn_long(3497);
	dataBufferOut_long( 102) <= dataBufferIn_long(3498);
	dataBufferOut_long( 845) <= dataBufferIn_long(3499);
	dataBufferOut_long(1588) <= dataBufferIn_long(3500);
	dataBufferOut_long(2331) <= dataBufferIn_long(3501);
	dataBufferOut_long(3074) <= dataBufferIn_long(3502);
	dataBufferOut_long(3817) <= dataBufferIn_long(3503);
	dataBufferOut_long(4560) <= dataBufferIn_long(3504);
	dataBufferOut_long(5303) <= dataBufferIn_long(3505);
	dataBufferOut_long(6046) <= dataBufferIn_long(3506);
	dataBufferOut_long( 645) <= dataBufferIn_long(3507);
	dataBufferOut_long(1388) <= dataBufferIn_long(3508);
	dataBufferOut_long(2131) <= dataBufferIn_long(3509);
	dataBufferOut_long(2874) <= dataBufferIn_long(3510);
	dataBufferOut_long(3617) <= dataBufferIn_long(3511);
	dataBufferOut_long(4360) <= dataBufferIn_long(3512);
	dataBufferOut_long(5103) <= dataBufferIn_long(3513);
	dataBufferOut_long(5846) <= dataBufferIn_long(3514);
	dataBufferOut_long( 445) <= dataBufferIn_long(3515);
	dataBufferOut_long(1188) <= dataBufferIn_long(3516);
	dataBufferOut_long(1931) <= dataBufferIn_long(3517);
	dataBufferOut_long(2674) <= dataBufferIn_long(3518);
	dataBufferOut_long(3417) <= dataBufferIn_long(3519);
	dataBufferOut_long(4160) <= dataBufferIn_long(3520);
	dataBufferOut_long(4903) <= dataBufferIn_long(3521);
	dataBufferOut_long(5646) <= dataBufferIn_long(3522);
	dataBufferOut_long( 245) <= dataBufferIn_long(3523);
	dataBufferOut_long( 988) <= dataBufferIn_long(3524);
	dataBufferOut_long(1731) <= dataBufferIn_long(3525);
	dataBufferOut_long(2474) <= dataBufferIn_long(3526);
	dataBufferOut_long(3217) <= dataBufferIn_long(3527);
	dataBufferOut_long(3960) <= dataBufferIn_long(3528);
	dataBufferOut_long(4703) <= dataBufferIn_long(3529);
	dataBufferOut_long(5446) <= dataBufferIn_long(3530);
	dataBufferOut_long(  45) <= dataBufferIn_long(3531);
	dataBufferOut_long( 788) <= dataBufferIn_long(3532);
	dataBufferOut_long(1531) <= dataBufferIn_long(3533);
	dataBufferOut_long(2274) <= dataBufferIn_long(3534);
	dataBufferOut_long(3017) <= dataBufferIn_long(3535);
	dataBufferOut_long(3760) <= dataBufferIn_long(3536);
	dataBufferOut_long(4503) <= dataBufferIn_long(3537);
	dataBufferOut_long(5246) <= dataBufferIn_long(3538);
	dataBufferOut_long(5989) <= dataBufferIn_long(3539);
	dataBufferOut_long( 588) <= dataBufferIn_long(3540);
	dataBufferOut_long(1331) <= dataBufferIn_long(3541);
	dataBufferOut_long(2074) <= dataBufferIn_long(3542);
	dataBufferOut_long(2817) <= dataBufferIn_long(3543);
	dataBufferOut_long(3560) <= dataBufferIn_long(3544);
	dataBufferOut_long(4303) <= dataBufferIn_long(3545);
	dataBufferOut_long(5046) <= dataBufferIn_long(3546);
	dataBufferOut_long(5789) <= dataBufferIn_long(3547);
	dataBufferOut_long( 388) <= dataBufferIn_long(3548);
	dataBufferOut_long(1131) <= dataBufferIn_long(3549);
	dataBufferOut_long(1874) <= dataBufferIn_long(3550);
	dataBufferOut_long(2617) <= dataBufferIn_long(3551);
	dataBufferOut_long(3360) <= dataBufferIn_long(3552);
	dataBufferOut_long(4103) <= dataBufferIn_long(3553);
	dataBufferOut_long(4846) <= dataBufferIn_long(3554);
	dataBufferOut_long(5589) <= dataBufferIn_long(3555);
	dataBufferOut_long( 188) <= dataBufferIn_long(3556);
	dataBufferOut_long( 931) <= dataBufferIn_long(3557);
	dataBufferOut_long(1674) <= dataBufferIn_long(3558);
	dataBufferOut_long(2417) <= dataBufferIn_long(3559);
	dataBufferOut_long(3160) <= dataBufferIn_long(3560);
	dataBufferOut_long(3903) <= dataBufferIn_long(3561);
	dataBufferOut_long(4646) <= dataBufferIn_long(3562);
	dataBufferOut_long(5389) <= dataBufferIn_long(3563);
	dataBufferOut_long(6132) <= dataBufferIn_long(3564);
	dataBufferOut_long( 731) <= dataBufferIn_long(3565);
	dataBufferOut_long(1474) <= dataBufferIn_long(3566);
	dataBufferOut_long(2217) <= dataBufferIn_long(3567);
	dataBufferOut_long(2960) <= dataBufferIn_long(3568);
	dataBufferOut_long(3703) <= dataBufferIn_long(3569);
	dataBufferOut_long(4446) <= dataBufferIn_long(3570);
	dataBufferOut_long(5189) <= dataBufferIn_long(3571);
	dataBufferOut_long(5932) <= dataBufferIn_long(3572);
	dataBufferOut_long( 531) <= dataBufferIn_long(3573);
	dataBufferOut_long(1274) <= dataBufferIn_long(3574);
	dataBufferOut_long(2017) <= dataBufferIn_long(3575);
	dataBufferOut_long(2760) <= dataBufferIn_long(3576);
	dataBufferOut_long(3503) <= dataBufferIn_long(3577);
	dataBufferOut_long(4246) <= dataBufferIn_long(3578);
	dataBufferOut_long(4989) <= dataBufferIn_long(3579);
	dataBufferOut_long(5732) <= dataBufferIn_long(3580);
	dataBufferOut_long( 331) <= dataBufferIn_long(3581);
	dataBufferOut_long(1074) <= dataBufferIn_long(3582);
	dataBufferOut_long(1817) <= dataBufferIn_long(3583);
	dataBufferOut_long(2560) <= dataBufferIn_long(3584);
	dataBufferOut_long(3303) <= dataBufferIn_long(3585);
	dataBufferOut_long(4046) <= dataBufferIn_long(3586);
	dataBufferOut_long(4789) <= dataBufferIn_long(3587);
	dataBufferOut_long(5532) <= dataBufferIn_long(3588);
	dataBufferOut_long( 131) <= dataBufferIn_long(3589);
	dataBufferOut_long( 874) <= dataBufferIn_long(3590);
	dataBufferOut_long(1617) <= dataBufferIn_long(3591);
	dataBufferOut_long(2360) <= dataBufferIn_long(3592);
	dataBufferOut_long(3103) <= dataBufferIn_long(3593);
	dataBufferOut_long(3846) <= dataBufferIn_long(3594);
	dataBufferOut_long(4589) <= dataBufferIn_long(3595);
	dataBufferOut_long(5332) <= dataBufferIn_long(3596);
	dataBufferOut_long(6075) <= dataBufferIn_long(3597);
	dataBufferOut_long( 674) <= dataBufferIn_long(3598);
	dataBufferOut_long(1417) <= dataBufferIn_long(3599);
	dataBufferOut_long(2160) <= dataBufferIn_long(3600);
	dataBufferOut_long(2903) <= dataBufferIn_long(3601);
	dataBufferOut_long(3646) <= dataBufferIn_long(3602);
	dataBufferOut_long(4389) <= dataBufferIn_long(3603);
	dataBufferOut_long(5132) <= dataBufferIn_long(3604);
	dataBufferOut_long(5875) <= dataBufferIn_long(3605);
	dataBufferOut_long( 474) <= dataBufferIn_long(3606);
	dataBufferOut_long(1217) <= dataBufferIn_long(3607);
	dataBufferOut_long(1960) <= dataBufferIn_long(3608);
	dataBufferOut_long(2703) <= dataBufferIn_long(3609);
	dataBufferOut_long(3446) <= dataBufferIn_long(3610);
	dataBufferOut_long(4189) <= dataBufferIn_long(3611);
	dataBufferOut_long(4932) <= dataBufferIn_long(3612);
	dataBufferOut_long(5675) <= dataBufferIn_long(3613);
	dataBufferOut_long( 274) <= dataBufferIn_long(3614);
	dataBufferOut_long(1017) <= dataBufferIn_long(3615);
	dataBufferOut_long(1760) <= dataBufferIn_long(3616);
	dataBufferOut_long(2503) <= dataBufferIn_long(3617);
	dataBufferOut_long(3246) <= dataBufferIn_long(3618);
	dataBufferOut_long(3989) <= dataBufferIn_long(3619);
	dataBufferOut_long(4732) <= dataBufferIn_long(3620);
	dataBufferOut_long(5475) <= dataBufferIn_long(3621);
	dataBufferOut_long(  74) <= dataBufferIn_long(3622);
	dataBufferOut_long( 817) <= dataBufferIn_long(3623);
	dataBufferOut_long(1560) <= dataBufferIn_long(3624);
	dataBufferOut_long(2303) <= dataBufferIn_long(3625);
	dataBufferOut_long(3046) <= dataBufferIn_long(3626);
	dataBufferOut_long(3789) <= dataBufferIn_long(3627);
	dataBufferOut_long(4532) <= dataBufferIn_long(3628);
	dataBufferOut_long(5275) <= dataBufferIn_long(3629);
	dataBufferOut_long(6018) <= dataBufferIn_long(3630);
	dataBufferOut_long( 617) <= dataBufferIn_long(3631);
	dataBufferOut_long(1360) <= dataBufferIn_long(3632);
	dataBufferOut_long(2103) <= dataBufferIn_long(3633);
	dataBufferOut_long(2846) <= dataBufferIn_long(3634);
	dataBufferOut_long(3589) <= dataBufferIn_long(3635);
	dataBufferOut_long(4332) <= dataBufferIn_long(3636);
	dataBufferOut_long(5075) <= dataBufferIn_long(3637);
	dataBufferOut_long(5818) <= dataBufferIn_long(3638);
	dataBufferOut_long( 417) <= dataBufferIn_long(3639);
	dataBufferOut_long(1160) <= dataBufferIn_long(3640);
	dataBufferOut_long(1903) <= dataBufferIn_long(3641);
	dataBufferOut_long(2646) <= dataBufferIn_long(3642);
	dataBufferOut_long(3389) <= dataBufferIn_long(3643);
	dataBufferOut_long(4132) <= dataBufferIn_long(3644);
	dataBufferOut_long(4875) <= dataBufferIn_long(3645);
	dataBufferOut_long(5618) <= dataBufferIn_long(3646);
	dataBufferOut_long( 217) <= dataBufferIn_long(3647);
	dataBufferOut_long( 960) <= dataBufferIn_long(3648);
	dataBufferOut_long(1703) <= dataBufferIn_long(3649);
	dataBufferOut_long(2446) <= dataBufferIn_long(3650);
	dataBufferOut_long(3189) <= dataBufferIn_long(3651);
	dataBufferOut_long(3932) <= dataBufferIn_long(3652);
	dataBufferOut_long(4675) <= dataBufferIn_long(3653);
	dataBufferOut_long(5418) <= dataBufferIn_long(3654);
	dataBufferOut_long(  17) <= dataBufferIn_long(3655);
	dataBufferOut_long( 760) <= dataBufferIn_long(3656);
	dataBufferOut_long(1503) <= dataBufferIn_long(3657);
	dataBufferOut_long(2246) <= dataBufferIn_long(3658);
	dataBufferOut_long(2989) <= dataBufferIn_long(3659);
	dataBufferOut_long(3732) <= dataBufferIn_long(3660);
	dataBufferOut_long(4475) <= dataBufferIn_long(3661);
	dataBufferOut_long(5218) <= dataBufferIn_long(3662);
	dataBufferOut_long(5961) <= dataBufferIn_long(3663);
	dataBufferOut_long( 560) <= dataBufferIn_long(3664);
	dataBufferOut_long(1303) <= dataBufferIn_long(3665);
	dataBufferOut_long(2046) <= dataBufferIn_long(3666);
	dataBufferOut_long(2789) <= dataBufferIn_long(3667);
	dataBufferOut_long(3532) <= dataBufferIn_long(3668);
	dataBufferOut_long(4275) <= dataBufferIn_long(3669);
	dataBufferOut_long(5018) <= dataBufferIn_long(3670);
	dataBufferOut_long(5761) <= dataBufferIn_long(3671);
	dataBufferOut_long( 360) <= dataBufferIn_long(3672);
	dataBufferOut_long(1103) <= dataBufferIn_long(3673);
	dataBufferOut_long(1846) <= dataBufferIn_long(3674);
	dataBufferOut_long(2589) <= dataBufferIn_long(3675);
	dataBufferOut_long(3332) <= dataBufferIn_long(3676);
	dataBufferOut_long(4075) <= dataBufferIn_long(3677);
	dataBufferOut_long(4818) <= dataBufferIn_long(3678);
	dataBufferOut_long(5561) <= dataBufferIn_long(3679);
	dataBufferOut_long( 160) <= dataBufferIn_long(3680);
	dataBufferOut_long( 903) <= dataBufferIn_long(3681);
	dataBufferOut_long(1646) <= dataBufferIn_long(3682);
	dataBufferOut_long(2389) <= dataBufferIn_long(3683);
	dataBufferOut_long(3132) <= dataBufferIn_long(3684);
	dataBufferOut_long(3875) <= dataBufferIn_long(3685);
	dataBufferOut_long(4618) <= dataBufferIn_long(3686);
	dataBufferOut_long(5361) <= dataBufferIn_long(3687);
	dataBufferOut_long(6104) <= dataBufferIn_long(3688);
	dataBufferOut_long( 703) <= dataBufferIn_long(3689);
	dataBufferOut_long(1446) <= dataBufferIn_long(3690);
	dataBufferOut_long(2189) <= dataBufferIn_long(3691);
	dataBufferOut_long(2932) <= dataBufferIn_long(3692);
	dataBufferOut_long(3675) <= dataBufferIn_long(3693);
	dataBufferOut_long(4418) <= dataBufferIn_long(3694);
	dataBufferOut_long(5161) <= dataBufferIn_long(3695);
	dataBufferOut_long(5904) <= dataBufferIn_long(3696);
	dataBufferOut_long( 503) <= dataBufferIn_long(3697);
	dataBufferOut_long(1246) <= dataBufferIn_long(3698);
	dataBufferOut_long(1989) <= dataBufferIn_long(3699);
	dataBufferOut_long(2732) <= dataBufferIn_long(3700);
	dataBufferOut_long(3475) <= dataBufferIn_long(3701);
	dataBufferOut_long(4218) <= dataBufferIn_long(3702);
	dataBufferOut_long(4961) <= dataBufferIn_long(3703);
	dataBufferOut_long(5704) <= dataBufferIn_long(3704);
	dataBufferOut_long( 303) <= dataBufferIn_long(3705);
	dataBufferOut_long(1046) <= dataBufferIn_long(3706);
	dataBufferOut_long(1789) <= dataBufferIn_long(3707);
	dataBufferOut_long(2532) <= dataBufferIn_long(3708);
	dataBufferOut_long(3275) <= dataBufferIn_long(3709);
	dataBufferOut_long(4018) <= dataBufferIn_long(3710);
	dataBufferOut_long(4761) <= dataBufferIn_long(3711);
	dataBufferOut_long(5504) <= dataBufferIn_long(3712);
	dataBufferOut_long( 103) <= dataBufferIn_long(3713);
	dataBufferOut_long( 846) <= dataBufferIn_long(3714);
	dataBufferOut_long(1589) <= dataBufferIn_long(3715);
	dataBufferOut_long(2332) <= dataBufferIn_long(3716);
	dataBufferOut_long(3075) <= dataBufferIn_long(3717);
	dataBufferOut_long(3818) <= dataBufferIn_long(3718);
	dataBufferOut_long(4561) <= dataBufferIn_long(3719);
	dataBufferOut_long(5304) <= dataBufferIn_long(3720);
	dataBufferOut_long(6047) <= dataBufferIn_long(3721);
	dataBufferOut_long( 646) <= dataBufferIn_long(3722);
	dataBufferOut_long(1389) <= dataBufferIn_long(3723);
	dataBufferOut_long(2132) <= dataBufferIn_long(3724);
	dataBufferOut_long(2875) <= dataBufferIn_long(3725);
	dataBufferOut_long(3618) <= dataBufferIn_long(3726);
	dataBufferOut_long(4361) <= dataBufferIn_long(3727);
	dataBufferOut_long(5104) <= dataBufferIn_long(3728);
	dataBufferOut_long(5847) <= dataBufferIn_long(3729);
	dataBufferOut_long( 446) <= dataBufferIn_long(3730);
	dataBufferOut_long(1189) <= dataBufferIn_long(3731);
	dataBufferOut_long(1932) <= dataBufferIn_long(3732);
	dataBufferOut_long(2675) <= dataBufferIn_long(3733);
	dataBufferOut_long(3418) <= dataBufferIn_long(3734);
	dataBufferOut_long(4161) <= dataBufferIn_long(3735);
	dataBufferOut_long(4904) <= dataBufferIn_long(3736);
	dataBufferOut_long(5647) <= dataBufferIn_long(3737);
	dataBufferOut_long( 246) <= dataBufferIn_long(3738);
	dataBufferOut_long( 989) <= dataBufferIn_long(3739);
	dataBufferOut_long(1732) <= dataBufferIn_long(3740);
	dataBufferOut_long(2475) <= dataBufferIn_long(3741);
	dataBufferOut_long(3218) <= dataBufferIn_long(3742);
	dataBufferOut_long(3961) <= dataBufferIn_long(3743);
	dataBufferOut_long(4704) <= dataBufferIn_long(3744);
	dataBufferOut_long(5447) <= dataBufferIn_long(3745);
	dataBufferOut_long(  46) <= dataBufferIn_long(3746);
	dataBufferOut_long( 789) <= dataBufferIn_long(3747);
	dataBufferOut_long(1532) <= dataBufferIn_long(3748);
	dataBufferOut_long(2275) <= dataBufferIn_long(3749);
	dataBufferOut_long(3018) <= dataBufferIn_long(3750);
	dataBufferOut_long(3761) <= dataBufferIn_long(3751);
	dataBufferOut_long(4504) <= dataBufferIn_long(3752);
	dataBufferOut_long(5247) <= dataBufferIn_long(3753);
	dataBufferOut_long(5990) <= dataBufferIn_long(3754);
	dataBufferOut_long( 589) <= dataBufferIn_long(3755);
	dataBufferOut_long(1332) <= dataBufferIn_long(3756);
	dataBufferOut_long(2075) <= dataBufferIn_long(3757);
	dataBufferOut_long(2818) <= dataBufferIn_long(3758);
	dataBufferOut_long(3561) <= dataBufferIn_long(3759);
	dataBufferOut_long(4304) <= dataBufferIn_long(3760);
	dataBufferOut_long(5047) <= dataBufferIn_long(3761);
	dataBufferOut_long(5790) <= dataBufferIn_long(3762);
	dataBufferOut_long( 389) <= dataBufferIn_long(3763);
	dataBufferOut_long(1132) <= dataBufferIn_long(3764);
	dataBufferOut_long(1875) <= dataBufferIn_long(3765);
	dataBufferOut_long(2618) <= dataBufferIn_long(3766);
	dataBufferOut_long(3361) <= dataBufferIn_long(3767);
	dataBufferOut_long(4104) <= dataBufferIn_long(3768);
	dataBufferOut_long(4847) <= dataBufferIn_long(3769);
	dataBufferOut_long(5590) <= dataBufferIn_long(3770);
	dataBufferOut_long( 189) <= dataBufferIn_long(3771);
	dataBufferOut_long( 932) <= dataBufferIn_long(3772);
	dataBufferOut_long(1675) <= dataBufferIn_long(3773);
	dataBufferOut_long(2418) <= dataBufferIn_long(3774);
	dataBufferOut_long(3161) <= dataBufferIn_long(3775);
	dataBufferOut_long(3904) <= dataBufferIn_long(3776);
	dataBufferOut_long(4647) <= dataBufferIn_long(3777);
	dataBufferOut_long(5390) <= dataBufferIn_long(3778);
	dataBufferOut_long(6133) <= dataBufferIn_long(3779);
	dataBufferOut_long( 732) <= dataBufferIn_long(3780);
	dataBufferOut_long(1475) <= dataBufferIn_long(3781);
	dataBufferOut_long(2218) <= dataBufferIn_long(3782);
	dataBufferOut_long(2961) <= dataBufferIn_long(3783);
	dataBufferOut_long(3704) <= dataBufferIn_long(3784);
	dataBufferOut_long(4447) <= dataBufferIn_long(3785);
	dataBufferOut_long(5190) <= dataBufferIn_long(3786);
	dataBufferOut_long(5933) <= dataBufferIn_long(3787);
	dataBufferOut_long( 532) <= dataBufferIn_long(3788);
	dataBufferOut_long(1275) <= dataBufferIn_long(3789);
	dataBufferOut_long(2018) <= dataBufferIn_long(3790);
	dataBufferOut_long(2761) <= dataBufferIn_long(3791);
	dataBufferOut_long(3504) <= dataBufferIn_long(3792);
	dataBufferOut_long(4247) <= dataBufferIn_long(3793);
	dataBufferOut_long(4990) <= dataBufferIn_long(3794);
	dataBufferOut_long(5733) <= dataBufferIn_long(3795);
	dataBufferOut_long( 332) <= dataBufferIn_long(3796);
	dataBufferOut_long(1075) <= dataBufferIn_long(3797);
	dataBufferOut_long(1818) <= dataBufferIn_long(3798);
	dataBufferOut_long(2561) <= dataBufferIn_long(3799);
	dataBufferOut_long(3304) <= dataBufferIn_long(3800);
	dataBufferOut_long(4047) <= dataBufferIn_long(3801);
	dataBufferOut_long(4790) <= dataBufferIn_long(3802);
	dataBufferOut_long(5533) <= dataBufferIn_long(3803);
	dataBufferOut_long( 132) <= dataBufferIn_long(3804);
	dataBufferOut_long( 875) <= dataBufferIn_long(3805);
	dataBufferOut_long(1618) <= dataBufferIn_long(3806);
	dataBufferOut_long(2361) <= dataBufferIn_long(3807);
	dataBufferOut_long(3104) <= dataBufferIn_long(3808);
	dataBufferOut_long(3847) <= dataBufferIn_long(3809);
	dataBufferOut_long(4590) <= dataBufferIn_long(3810);
	dataBufferOut_long(5333) <= dataBufferIn_long(3811);
	dataBufferOut_long(6076) <= dataBufferIn_long(3812);
	dataBufferOut_long( 675) <= dataBufferIn_long(3813);
	dataBufferOut_long(1418) <= dataBufferIn_long(3814);
	dataBufferOut_long(2161) <= dataBufferIn_long(3815);
	dataBufferOut_long(2904) <= dataBufferIn_long(3816);
	dataBufferOut_long(3647) <= dataBufferIn_long(3817);
	dataBufferOut_long(4390) <= dataBufferIn_long(3818);
	dataBufferOut_long(5133) <= dataBufferIn_long(3819);
	dataBufferOut_long(5876) <= dataBufferIn_long(3820);
	dataBufferOut_long( 475) <= dataBufferIn_long(3821);
	dataBufferOut_long(1218) <= dataBufferIn_long(3822);
	dataBufferOut_long(1961) <= dataBufferIn_long(3823);
	dataBufferOut_long(2704) <= dataBufferIn_long(3824);
	dataBufferOut_long(3447) <= dataBufferIn_long(3825);
	dataBufferOut_long(4190) <= dataBufferIn_long(3826);
	dataBufferOut_long(4933) <= dataBufferIn_long(3827);
	dataBufferOut_long(5676) <= dataBufferIn_long(3828);
	dataBufferOut_long( 275) <= dataBufferIn_long(3829);
	dataBufferOut_long(1018) <= dataBufferIn_long(3830);
	dataBufferOut_long(1761) <= dataBufferIn_long(3831);
	dataBufferOut_long(2504) <= dataBufferIn_long(3832);
	dataBufferOut_long(3247) <= dataBufferIn_long(3833);
	dataBufferOut_long(3990) <= dataBufferIn_long(3834);
	dataBufferOut_long(4733) <= dataBufferIn_long(3835);
	dataBufferOut_long(5476) <= dataBufferIn_long(3836);
	dataBufferOut_long(  75) <= dataBufferIn_long(3837);
	dataBufferOut_long( 818) <= dataBufferIn_long(3838);
	dataBufferOut_long(1561) <= dataBufferIn_long(3839);
	dataBufferOut_long(2304) <= dataBufferIn_long(3840);
	dataBufferOut_long(3047) <= dataBufferIn_long(3841);
	dataBufferOut_long(3790) <= dataBufferIn_long(3842);
	dataBufferOut_long(4533) <= dataBufferIn_long(3843);
	dataBufferOut_long(5276) <= dataBufferIn_long(3844);
	dataBufferOut_long(6019) <= dataBufferIn_long(3845);
	dataBufferOut_long( 618) <= dataBufferIn_long(3846);
	dataBufferOut_long(1361) <= dataBufferIn_long(3847);
	dataBufferOut_long(2104) <= dataBufferIn_long(3848);
	dataBufferOut_long(2847) <= dataBufferIn_long(3849);
	dataBufferOut_long(3590) <= dataBufferIn_long(3850);
	dataBufferOut_long(4333) <= dataBufferIn_long(3851);
	dataBufferOut_long(5076) <= dataBufferIn_long(3852);
	dataBufferOut_long(5819) <= dataBufferIn_long(3853);
	dataBufferOut_long( 418) <= dataBufferIn_long(3854);
	dataBufferOut_long(1161) <= dataBufferIn_long(3855);
	dataBufferOut_long(1904) <= dataBufferIn_long(3856);
	dataBufferOut_long(2647) <= dataBufferIn_long(3857);
	dataBufferOut_long(3390) <= dataBufferIn_long(3858);
	dataBufferOut_long(4133) <= dataBufferIn_long(3859);
	dataBufferOut_long(4876) <= dataBufferIn_long(3860);
	dataBufferOut_long(5619) <= dataBufferIn_long(3861);
	dataBufferOut_long( 218) <= dataBufferIn_long(3862);
	dataBufferOut_long( 961) <= dataBufferIn_long(3863);
	dataBufferOut_long(1704) <= dataBufferIn_long(3864);
	dataBufferOut_long(2447) <= dataBufferIn_long(3865);
	dataBufferOut_long(3190) <= dataBufferIn_long(3866);
	dataBufferOut_long(3933) <= dataBufferIn_long(3867);
	dataBufferOut_long(4676) <= dataBufferIn_long(3868);
	dataBufferOut_long(5419) <= dataBufferIn_long(3869);
	dataBufferOut_long(  18) <= dataBufferIn_long(3870);
	dataBufferOut_long( 761) <= dataBufferIn_long(3871);
	dataBufferOut_long(1504) <= dataBufferIn_long(3872);
	dataBufferOut_long(2247) <= dataBufferIn_long(3873);
	dataBufferOut_long(2990) <= dataBufferIn_long(3874);
	dataBufferOut_long(3733) <= dataBufferIn_long(3875);
	dataBufferOut_long(4476) <= dataBufferIn_long(3876);
	dataBufferOut_long(5219) <= dataBufferIn_long(3877);
	dataBufferOut_long(5962) <= dataBufferIn_long(3878);
	dataBufferOut_long( 561) <= dataBufferIn_long(3879);
	dataBufferOut_long(1304) <= dataBufferIn_long(3880);
	dataBufferOut_long(2047) <= dataBufferIn_long(3881);
	dataBufferOut_long(2790) <= dataBufferIn_long(3882);
	dataBufferOut_long(3533) <= dataBufferIn_long(3883);
	dataBufferOut_long(4276) <= dataBufferIn_long(3884);
	dataBufferOut_long(5019) <= dataBufferIn_long(3885);
	dataBufferOut_long(5762) <= dataBufferIn_long(3886);
	dataBufferOut_long( 361) <= dataBufferIn_long(3887);
	dataBufferOut_long(1104) <= dataBufferIn_long(3888);
	dataBufferOut_long(1847) <= dataBufferIn_long(3889);
	dataBufferOut_long(2590) <= dataBufferIn_long(3890);
	dataBufferOut_long(3333) <= dataBufferIn_long(3891);
	dataBufferOut_long(4076) <= dataBufferIn_long(3892);
	dataBufferOut_long(4819) <= dataBufferIn_long(3893);
	dataBufferOut_long(5562) <= dataBufferIn_long(3894);
	dataBufferOut_long( 161) <= dataBufferIn_long(3895);
	dataBufferOut_long( 904) <= dataBufferIn_long(3896);
	dataBufferOut_long(1647) <= dataBufferIn_long(3897);
	dataBufferOut_long(2390) <= dataBufferIn_long(3898);
	dataBufferOut_long(3133) <= dataBufferIn_long(3899);
	dataBufferOut_long(3876) <= dataBufferIn_long(3900);
	dataBufferOut_long(4619) <= dataBufferIn_long(3901);
	dataBufferOut_long(5362) <= dataBufferIn_long(3902);
	dataBufferOut_long(6105) <= dataBufferIn_long(3903);
	dataBufferOut_long( 704) <= dataBufferIn_long(3904);
	dataBufferOut_long(1447) <= dataBufferIn_long(3905);
	dataBufferOut_long(2190) <= dataBufferIn_long(3906);
	dataBufferOut_long(2933) <= dataBufferIn_long(3907);
	dataBufferOut_long(3676) <= dataBufferIn_long(3908);
	dataBufferOut_long(4419) <= dataBufferIn_long(3909);
	dataBufferOut_long(5162) <= dataBufferIn_long(3910);
	dataBufferOut_long(5905) <= dataBufferIn_long(3911);
	dataBufferOut_long( 504) <= dataBufferIn_long(3912);
	dataBufferOut_long(1247) <= dataBufferIn_long(3913);
	dataBufferOut_long(1990) <= dataBufferIn_long(3914);
	dataBufferOut_long(2733) <= dataBufferIn_long(3915);
	dataBufferOut_long(3476) <= dataBufferIn_long(3916);
	dataBufferOut_long(4219) <= dataBufferIn_long(3917);
	dataBufferOut_long(4962) <= dataBufferIn_long(3918);
	dataBufferOut_long(5705) <= dataBufferIn_long(3919);
	dataBufferOut_long( 304) <= dataBufferIn_long(3920);
	dataBufferOut_long(1047) <= dataBufferIn_long(3921);
	dataBufferOut_long(1790) <= dataBufferIn_long(3922);
	dataBufferOut_long(2533) <= dataBufferIn_long(3923);
	dataBufferOut_long(3276) <= dataBufferIn_long(3924);
	dataBufferOut_long(4019) <= dataBufferIn_long(3925);
	dataBufferOut_long(4762) <= dataBufferIn_long(3926);
	dataBufferOut_long(5505) <= dataBufferIn_long(3927);
	dataBufferOut_long( 104) <= dataBufferIn_long(3928);
	dataBufferOut_long( 847) <= dataBufferIn_long(3929);
	dataBufferOut_long(1590) <= dataBufferIn_long(3930);
	dataBufferOut_long(2333) <= dataBufferIn_long(3931);
	dataBufferOut_long(3076) <= dataBufferIn_long(3932);
	dataBufferOut_long(3819) <= dataBufferIn_long(3933);
	dataBufferOut_long(4562) <= dataBufferIn_long(3934);
	dataBufferOut_long(5305) <= dataBufferIn_long(3935);
	dataBufferOut_long(6048) <= dataBufferIn_long(3936);
	dataBufferOut_long( 647) <= dataBufferIn_long(3937);
	dataBufferOut_long(1390) <= dataBufferIn_long(3938);
	dataBufferOut_long(2133) <= dataBufferIn_long(3939);
	dataBufferOut_long(2876) <= dataBufferIn_long(3940);
	dataBufferOut_long(3619) <= dataBufferIn_long(3941);
	dataBufferOut_long(4362) <= dataBufferIn_long(3942);
	dataBufferOut_long(5105) <= dataBufferIn_long(3943);
	dataBufferOut_long(5848) <= dataBufferIn_long(3944);
	dataBufferOut_long( 447) <= dataBufferIn_long(3945);
	dataBufferOut_long(1190) <= dataBufferIn_long(3946);
	dataBufferOut_long(1933) <= dataBufferIn_long(3947);
	dataBufferOut_long(2676) <= dataBufferIn_long(3948);
	dataBufferOut_long(3419) <= dataBufferIn_long(3949);
	dataBufferOut_long(4162) <= dataBufferIn_long(3950);
	dataBufferOut_long(4905) <= dataBufferIn_long(3951);
	dataBufferOut_long(5648) <= dataBufferIn_long(3952);
	dataBufferOut_long( 247) <= dataBufferIn_long(3953);
	dataBufferOut_long( 990) <= dataBufferIn_long(3954);
	dataBufferOut_long(1733) <= dataBufferIn_long(3955);
	dataBufferOut_long(2476) <= dataBufferIn_long(3956);
	dataBufferOut_long(3219) <= dataBufferIn_long(3957);
	dataBufferOut_long(3962) <= dataBufferIn_long(3958);
	dataBufferOut_long(4705) <= dataBufferIn_long(3959);
	dataBufferOut_long(5448) <= dataBufferIn_long(3960);
	dataBufferOut_long(  47) <= dataBufferIn_long(3961);
	dataBufferOut_long( 790) <= dataBufferIn_long(3962);
	dataBufferOut_long(1533) <= dataBufferIn_long(3963);
	dataBufferOut_long(2276) <= dataBufferIn_long(3964);
	dataBufferOut_long(3019) <= dataBufferIn_long(3965);
	dataBufferOut_long(3762) <= dataBufferIn_long(3966);
	dataBufferOut_long(4505) <= dataBufferIn_long(3967);
	dataBufferOut_long(5248) <= dataBufferIn_long(3968);
	dataBufferOut_long(5991) <= dataBufferIn_long(3969);
	dataBufferOut_long( 590) <= dataBufferIn_long(3970);
	dataBufferOut_long(1333) <= dataBufferIn_long(3971);
	dataBufferOut_long(2076) <= dataBufferIn_long(3972);
	dataBufferOut_long(2819) <= dataBufferIn_long(3973);
	dataBufferOut_long(3562) <= dataBufferIn_long(3974);
	dataBufferOut_long(4305) <= dataBufferIn_long(3975);
	dataBufferOut_long(5048) <= dataBufferIn_long(3976);
	dataBufferOut_long(5791) <= dataBufferIn_long(3977);
	dataBufferOut_long( 390) <= dataBufferIn_long(3978);
	dataBufferOut_long(1133) <= dataBufferIn_long(3979);
	dataBufferOut_long(1876) <= dataBufferIn_long(3980);
	dataBufferOut_long(2619) <= dataBufferIn_long(3981);
	dataBufferOut_long(3362) <= dataBufferIn_long(3982);
	dataBufferOut_long(4105) <= dataBufferIn_long(3983);
	dataBufferOut_long(4848) <= dataBufferIn_long(3984);
	dataBufferOut_long(5591) <= dataBufferIn_long(3985);
	dataBufferOut_long( 190) <= dataBufferIn_long(3986);
	dataBufferOut_long( 933) <= dataBufferIn_long(3987);
	dataBufferOut_long(1676) <= dataBufferIn_long(3988);
	dataBufferOut_long(2419) <= dataBufferIn_long(3989);
	dataBufferOut_long(3162) <= dataBufferIn_long(3990);
	dataBufferOut_long(3905) <= dataBufferIn_long(3991);
	dataBufferOut_long(4648) <= dataBufferIn_long(3992);
	dataBufferOut_long(5391) <= dataBufferIn_long(3993);
	dataBufferOut_long(6134) <= dataBufferIn_long(3994);
	dataBufferOut_long( 733) <= dataBufferIn_long(3995);
	dataBufferOut_long(1476) <= dataBufferIn_long(3996);
	dataBufferOut_long(2219) <= dataBufferIn_long(3997);
	dataBufferOut_long(2962) <= dataBufferIn_long(3998);
	dataBufferOut_long(3705) <= dataBufferIn_long(3999);
	dataBufferOut_long(4448) <= dataBufferIn_long(4000);
	dataBufferOut_long(5191) <= dataBufferIn_long(4001);
	dataBufferOut_long(5934) <= dataBufferIn_long(4002);
	dataBufferOut_long( 533) <= dataBufferIn_long(4003);
	dataBufferOut_long(1276) <= dataBufferIn_long(4004);
	dataBufferOut_long(2019) <= dataBufferIn_long(4005);
	dataBufferOut_long(2762) <= dataBufferIn_long(4006);
	dataBufferOut_long(3505) <= dataBufferIn_long(4007);
	dataBufferOut_long(4248) <= dataBufferIn_long(4008);
	dataBufferOut_long(4991) <= dataBufferIn_long(4009);
	dataBufferOut_long(5734) <= dataBufferIn_long(4010);
	dataBufferOut_long( 333) <= dataBufferIn_long(4011);
	dataBufferOut_long(1076) <= dataBufferIn_long(4012);
	dataBufferOut_long(1819) <= dataBufferIn_long(4013);
	dataBufferOut_long(2562) <= dataBufferIn_long(4014);
	dataBufferOut_long(3305) <= dataBufferIn_long(4015);
	dataBufferOut_long(4048) <= dataBufferIn_long(4016);
	dataBufferOut_long(4791) <= dataBufferIn_long(4017);
	dataBufferOut_long(5534) <= dataBufferIn_long(4018);
	dataBufferOut_long( 133) <= dataBufferIn_long(4019);
	dataBufferOut_long( 876) <= dataBufferIn_long(4020);
	dataBufferOut_long(1619) <= dataBufferIn_long(4021);
	dataBufferOut_long(2362) <= dataBufferIn_long(4022);
	dataBufferOut_long(3105) <= dataBufferIn_long(4023);
	dataBufferOut_long(3848) <= dataBufferIn_long(4024);
	dataBufferOut_long(4591) <= dataBufferIn_long(4025);
	dataBufferOut_long(5334) <= dataBufferIn_long(4026);
	dataBufferOut_long(6077) <= dataBufferIn_long(4027);
	dataBufferOut_long( 676) <= dataBufferIn_long(4028);
	dataBufferOut_long(1419) <= dataBufferIn_long(4029);
	dataBufferOut_long(2162) <= dataBufferIn_long(4030);
	dataBufferOut_long(2905) <= dataBufferIn_long(4031);
	dataBufferOut_long(3648) <= dataBufferIn_long(4032);
	dataBufferOut_long(4391) <= dataBufferIn_long(4033);
	dataBufferOut_long(5134) <= dataBufferIn_long(4034);
	dataBufferOut_long(5877) <= dataBufferIn_long(4035);
	dataBufferOut_long( 476) <= dataBufferIn_long(4036);
	dataBufferOut_long(1219) <= dataBufferIn_long(4037);
	dataBufferOut_long(1962) <= dataBufferIn_long(4038);
	dataBufferOut_long(2705) <= dataBufferIn_long(4039);
	dataBufferOut_long(3448) <= dataBufferIn_long(4040);
	dataBufferOut_long(4191) <= dataBufferIn_long(4041);
	dataBufferOut_long(4934) <= dataBufferIn_long(4042);
	dataBufferOut_long(5677) <= dataBufferIn_long(4043);
	dataBufferOut_long( 276) <= dataBufferIn_long(4044);
	dataBufferOut_long(1019) <= dataBufferIn_long(4045);
	dataBufferOut_long(1762) <= dataBufferIn_long(4046);
	dataBufferOut_long(2505) <= dataBufferIn_long(4047);
	dataBufferOut_long(3248) <= dataBufferIn_long(4048);
	dataBufferOut_long(3991) <= dataBufferIn_long(4049);
	dataBufferOut_long(4734) <= dataBufferIn_long(4050);
	dataBufferOut_long(5477) <= dataBufferIn_long(4051);
	dataBufferOut_long(  76) <= dataBufferIn_long(4052);
	dataBufferOut_long( 819) <= dataBufferIn_long(4053);
	dataBufferOut_long(1562) <= dataBufferIn_long(4054);
	dataBufferOut_long(2305) <= dataBufferIn_long(4055);
	dataBufferOut_long(3048) <= dataBufferIn_long(4056);
	dataBufferOut_long(3791) <= dataBufferIn_long(4057);
	dataBufferOut_long(4534) <= dataBufferIn_long(4058);
	dataBufferOut_long(5277) <= dataBufferIn_long(4059);
	dataBufferOut_long(6020) <= dataBufferIn_long(4060);
	dataBufferOut_long( 619) <= dataBufferIn_long(4061);
	dataBufferOut_long(1362) <= dataBufferIn_long(4062);
	dataBufferOut_long(2105) <= dataBufferIn_long(4063);
	dataBufferOut_long(2848) <= dataBufferIn_long(4064);
	dataBufferOut_long(3591) <= dataBufferIn_long(4065);
	dataBufferOut_long(4334) <= dataBufferIn_long(4066);
	dataBufferOut_long(5077) <= dataBufferIn_long(4067);
	dataBufferOut_long(5820) <= dataBufferIn_long(4068);
	dataBufferOut_long( 419) <= dataBufferIn_long(4069);
	dataBufferOut_long(1162) <= dataBufferIn_long(4070);
	dataBufferOut_long(1905) <= dataBufferIn_long(4071);
	dataBufferOut_long(2648) <= dataBufferIn_long(4072);
	dataBufferOut_long(3391) <= dataBufferIn_long(4073);
	dataBufferOut_long(4134) <= dataBufferIn_long(4074);
	dataBufferOut_long(4877) <= dataBufferIn_long(4075);
	dataBufferOut_long(5620) <= dataBufferIn_long(4076);
	dataBufferOut_long( 219) <= dataBufferIn_long(4077);
	dataBufferOut_long( 962) <= dataBufferIn_long(4078);
	dataBufferOut_long(1705) <= dataBufferIn_long(4079);
	dataBufferOut_long(2448) <= dataBufferIn_long(4080);
	dataBufferOut_long(3191) <= dataBufferIn_long(4081);
	dataBufferOut_long(3934) <= dataBufferIn_long(4082);
	dataBufferOut_long(4677) <= dataBufferIn_long(4083);
	dataBufferOut_long(5420) <= dataBufferIn_long(4084);
	dataBufferOut_long(  19) <= dataBufferIn_long(4085);
	dataBufferOut_long( 762) <= dataBufferIn_long(4086);
	dataBufferOut_long(1505) <= dataBufferIn_long(4087);
	dataBufferOut_long(2248) <= dataBufferIn_long(4088);
	dataBufferOut_long(2991) <= dataBufferIn_long(4089);
	dataBufferOut_long(3734) <= dataBufferIn_long(4090);
	dataBufferOut_long(4477) <= dataBufferIn_long(4091);
	dataBufferOut_long(5220) <= dataBufferIn_long(4092);
	dataBufferOut_long(5963) <= dataBufferIn_long(4093);
	dataBufferOut_long( 562) <= dataBufferIn_long(4094);
	dataBufferOut_long(1305) <= dataBufferIn_long(4095);
	dataBufferOut_long(2048) <= dataBufferIn_long(4096);
	dataBufferOut_long(2791) <= dataBufferIn_long(4097);
	dataBufferOut_long(3534) <= dataBufferIn_long(4098);
	dataBufferOut_long(4277) <= dataBufferIn_long(4099);
	dataBufferOut_long(5020) <= dataBufferIn_long(4100);
	dataBufferOut_long(5763) <= dataBufferIn_long(4101);
	dataBufferOut_long( 362) <= dataBufferIn_long(4102);
	dataBufferOut_long(1105) <= dataBufferIn_long(4103);
	dataBufferOut_long(1848) <= dataBufferIn_long(4104);
	dataBufferOut_long(2591) <= dataBufferIn_long(4105);
	dataBufferOut_long(3334) <= dataBufferIn_long(4106);
	dataBufferOut_long(4077) <= dataBufferIn_long(4107);
	dataBufferOut_long(4820) <= dataBufferIn_long(4108);
	dataBufferOut_long(5563) <= dataBufferIn_long(4109);
	dataBufferOut_long( 162) <= dataBufferIn_long(4110);
	dataBufferOut_long( 905) <= dataBufferIn_long(4111);
	dataBufferOut_long(1648) <= dataBufferIn_long(4112);
	dataBufferOut_long(2391) <= dataBufferIn_long(4113);
	dataBufferOut_long(3134) <= dataBufferIn_long(4114);
	dataBufferOut_long(3877) <= dataBufferIn_long(4115);
	dataBufferOut_long(4620) <= dataBufferIn_long(4116);
	dataBufferOut_long(5363) <= dataBufferIn_long(4117);
	dataBufferOut_long(6106) <= dataBufferIn_long(4118);
	dataBufferOut_long( 705) <= dataBufferIn_long(4119);
	dataBufferOut_long(1448) <= dataBufferIn_long(4120);
	dataBufferOut_long(2191) <= dataBufferIn_long(4121);
	dataBufferOut_long(2934) <= dataBufferIn_long(4122);
	dataBufferOut_long(3677) <= dataBufferIn_long(4123);
	dataBufferOut_long(4420) <= dataBufferIn_long(4124);
	dataBufferOut_long(5163) <= dataBufferIn_long(4125);
	dataBufferOut_long(5906) <= dataBufferIn_long(4126);
	dataBufferOut_long( 505) <= dataBufferIn_long(4127);
	dataBufferOut_long(1248) <= dataBufferIn_long(4128);
	dataBufferOut_long(1991) <= dataBufferIn_long(4129);
	dataBufferOut_long(2734) <= dataBufferIn_long(4130);
	dataBufferOut_long(3477) <= dataBufferIn_long(4131);
	dataBufferOut_long(4220) <= dataBufferIn_long(4132);
	dataBufferOut_long(4963) <= dataBufferIn_long(4133);
	dataBufferOut_long(5706) <= dataBufferIn_long(4134);
	dataBufferOut_long( 305) <= dataBufferIn_long(4135);
	dataBufferOut_long(1048) <= dataBufferIn_long(4136);
	dataBufferOut_long(1791) <= dataBufferIn_long(4137);
	dataBufferOut_long(2534) <= dataBufferIn_long(4138);
	dataBufferOut_long(3277) <= dataBufferIn_long(4139);
	dataBufferOut_long(4020) <= dataBufferIn_long(4140);
	dataBufferOut_long(4763) <= dataBufferIn_long(4141);
	dataBufferOut_long(5506) <= dataBufferIn_long(4142);
	dataBufferOut_long( 105) <= dataBufferIn_long(4143);
	dataBufferOut_long( 848) <= dataBufferIn_long(4144);
	dataBufferOut_long(1591) <= dataBufferIn_long(4145);
	dataBufferOut_long(2334) <= dataBufferIn_long(4146);
	dataBufferOut_long(3077) <= dataBufferIn_long(4147);
	dataBufferOut_long(3820) <= dataBufferIn_long(4148);
	dataBufferOut_long(4563) <= dataBufferIn_long(4149);
	dataBufferOut_long(5306) <= dataBufferIn_long(4150);
	dataBufferOut_long(6049) <= dataBufferIn_long(4151);
	dataBufferOut_long( 648) <= dataBufferIn_long(4152);
	dataBufferOut_long(1391) <= dataBufferIn_long(4153);
	dataBufferOut_long(2134) <= dataBufferIn_long(4154);
	dataBufferOut_long(2877) <= dataBufferIn_long(4155);
	dataBufferOut_long(3620) <= dataBufferIn_long(4156);
	dataBufferOut_long(4363) <= dataBufferIn_long(4157);
	dataBufferOut_long(5106) <= dataBufferIn_long(4158);
	dataBufferOut_long(5849) <= dataBufferIn_long(4159);
	dataBufferOut_long( 448) <= dataBufferIn_long(4160);
	dataBufferOut_long(1191) <= dataBufferIn_long(4161);
	dataBufferOut_long(1934) <= dataBufferIn_long(4162);
	dataBufferOut_long(2677) <= dataBufferIn_long(4163);
	dataBufferOut_long(3420) <= dataBufferIn_long(4164);
	dataBufferOut_long(4163) <= dataBufferIn_long(4165);
	dataBufferOut_long(4906) <= dataBufferIn_long(4166);
	dataBufferOut_long(5649) <= dataBufferIn_long(4167);
	dataBufferOut_long( 248) <= dataBufferIn_long(4168);
	dataBufferOut_long( 991) <= dataBufferIn_long(4169);
	dataBufferOut_long(1734) <= dataBufferIn_long(4170);
	dataBufferOut_long(2477) <= dataBufferIn_long(4171);
	dataBufferOut_long(3220) <= dataBufferIn_long(4172);
	dataBufferOut_long(3963) <= dataBufferIn_long(4173);
	dataBufferOut_long(4706) <= dataBufferIn_long(4174);
	dataBufferOut_long(5449) <= dataBufferIn_long(4175);
	dataBufferOut_long(  48) <= dataBufferIn_long(4176);
	dataBufferOut_long( 791) <= dataBufferIn_long(4177);
	dataBufferOut_long(1534) <= dataBufferIn_long(4178);
	dataBufferOut_long(2277) <= dataBufferIn_long(4179);
	dataBufferOut_long(3020) <= dataBufferIn_long(4180);
	dataBufferOut_long(3763) <= dataBufferIn_long(4181);
	dataBufferOut_long(4506) <= dataBufferIn_long(4182);
	dataBufferOut_long(5249) <= dataBufferIn_long(4183);
	dataBufferOut_long(5992) <= dataBufferIn_long(4184);
	dataBufferOut_long( 591) <= dataBufferIn_long(4185);
	dataBufferOut_long(1334) <= dataBufferIn_long(4186);
	dataBufferOut_long(2077) <= dataBufferIn_long(4187);
	dataBufferOut_long(2820) <= dataBufferIn_long(4188);
	dataBufferOut_long(3563) <= dataBufferIn_long(4189);
	dataBufferOut_long(4306) <= dataBufferIn_long(4190);
	dataBufferOut_long(5049) <= dataBufferIn_long(4191);
	dataBufferOut_long(5792) <= dataBufferIn_long(4192);
	dataBufferOut_long( 391) <= dataBufferIn_long(4193);
	dataBufferOut_long(1134) <= dataBufferIn_long(4194);
	dataBufferOut_long(1877) <= dataBufferIn_long(4195);
	dataBufferOut_long(2620) <= dataBufferIn_long(4196);
	dataBufferOut_long(3363) <= dataBufferIn_long(4197);
	dataBufferOut_long(4106) <= dataBufferIn_long(4198);
	dataBufferOut_long(4849) <= dataBufferIn_long(4199);
	dataBufferOut_long(5592) <= dataBufferIn_long(4200);
	dataBufferOut_long( 191) <= dataBufferIn_long(4201);
	dataBufferOut_long( 934) <= dataBufferIn_long(4202);
	dataBufferOut_long(1677) <= dataBufferIn_long(4203);
	dataBufferOut_long(2420) <= dataBufferIn_long(4204);
	dataBufferOut_long(3163) <= dataBufferIn_long(4205);
	dataBufferOut_long(3906) <= dataBufferIn_long(4206);
	dataBufferOut_long(4649) <= dataBufferIn_long(4207);
	dataBufferOut_long(5392) <= dataBufferIn_long(4208);
	dataBufferOut_long(6135) <= dataBufferIn_long(4209);
	dataBufferOut_long( 734) <= dataBufferIn_long(4210);
	dataBufferOut_long(1477) <= dataBufferIn_long(4211);
	dataBufferOut_long(2220) <= dataBufferIn_long(4212);
	dataBufferOut_long(2963) <= dataBufferIn_long(4213);
	dataBufferOut_long(3706) <= dataBufferIn_long(4214);
	dataBufferOut_long(4449) <= dataBufferIn_long(4215);
	dataBufferOut_long(5192) <= dataBufferIn_long(4216);
	dataBufferOut_long(5935) <= dataBufferIn_long(4217);
	dataBufferOut_long( 534) <= dataBufferIn_long(4218);
	dataBufferOut_long(1277) <= dataBufferIn_long(4219);
	dataBufferOut_long(2020) <= dataBufferIn_long(4220);
	dataBufferOut_long(2763) <= dataBufferIn_long(4221);
	dataBufferOut_long(3506) <= dataBufferIn_long(4222);
	dataBufferOut_long(4249) <= dataBufferIn_long(4223);
	dataBufferOut_long(4992) <= dataBufferIn_long(4224);
	dataBufferOut_long(5735) <= dataBufferIn_long(4225);
	dataBufferOut_long( 334) <= dataBufferIn_long(4226);
	dataBufferOut_long(1077) <= dataBufferIn_long(4227);
	dataBufferOut_long(1820) <= dataBufferIn_long(4228);
	dataBufferOut_long(2563) <= dataBufferIn_long(4229);
	dataBufferOut_long(3306) <= dataBufferIn_long(4230);
	dataBufferOut_long(4049) <= dataBufferIn_long(4231);
	dataBufferOut_long(4792) <= dataBufferIn_long(4232);
	dataBufferOut_long(5535) <= dataBufferIn_long(4233);
	dataBufferOut_long( 134) <= dataBufferIn_long(4234);
	dataBufferOut_long( 877) <= dataBufferIn_long(4235);
	dataBufferOut_long(1620) <= dataBufferIn_long(4236);
	dataBufferOut_long(2363) <= dataBufferIn_long(4237);
	dataBufferOut_long(3106) <= dataBufferIn_long(4238);
	dataBufferOut_long(3849) <= dataBufferIn_long(4239);
	dataBufferOut_long(4592) <= dataBufferIn_long(4240);
	dataBufferOut_long(5335) <= dataBufferIn_long(4241);
	dataBufferOut_long(6078) <= dataBufferIn_long(4242);
	dataBufferOut_long( 677) <= dataBufferIn_long(4243);
	dataBufferOut_long(1420) <= dataBufferIn_long(4244);
	dataBufferOut_long(2163) <= dataBufferIn_long(4245);
	dataBufferOut_long(2906) <= dataBufferIn_long(4246);
	dataBufferOut_long(3649) <= dataBufferIn_long(4247);
	dataBufferOut_long(4392) <= dataBufferIn_long(4248);
	dataBufferOut_long(5135) <= dataBufferIn_long(4249);
	dataBufferOut_long(5878) <= dataBufferIn_long(4250);
	dataBufferOut_long( 477) <= dataBufferIn_long(4251);
	dataBufferOut_long(1220) <= dataBufferIn_long(4252);
	dataBufferOut_long(1963) <= dataBufferIn_long(4253);
	dataBufferOut_long(2706) <= dataBufferIn_long(4254);
	dataBufferOut_long(3449) <= dataBufferIn_long(4255);
	dataBufferOut_long(4192) <= dataBufferIn_long(4256);
	dataBufferOut_long(4935) <= dataBufferIn_long(4257);
	dataBufferOut_long(5678) <= dataBufferIn_long(4258);
	dataBufferOut_long( 277) <= dataBufferIn_long(4259);
	dataBufferOut_long(1020) <= dataBufferIn_long(4260);
	dataBufferOut_long(1763) <= dataBufferIn_long(4261);
	dataBufferOut_long(2506) <= dataBufferIn_long(4262);
	dataBufferOut_long(3249) <= dataBufferIn_long(4263);
	dataBufferOut_long(3992) <= dataBufferIn_long(4264);
	dataBufferOut_long(4735) <= dataBufferIn_long(4265);
	dataBufferOut_long(5478) <= dataBufferIn_long(4266);
	dataBufferOut_long(  77) <= dataBufferIn_long(4267);
	dataBufferOut_long( 820) <= dataBufferIn_long(4268);
	dataBufferOut_long(1563) <= dataBufferIn_long(4269);
	dataBufferOut_long(2306) <= dataBufferIn_long(4270);
	dataBufferOut_long(3049) <= dataBufferIn_long(4271);
	dataBufferOut_long(3792) <= dataBufferIn_long(4272);
	dataBufferOut_long(4535) <= dataBufferIn_long(4273);
	dataBufferOut_long(5278) <= dataBufferIn_long(4274);
	dataBufferOut_long(6021) <= dataBufferIn_long(4275);
	dataBufferOut_long( 620) <= dataBufferIn_long(4276);
	dataBufferOut_long(1363) <= dataBufferIn_long(4277);
	dataBufferOut_long(2106) <= dataBufferIn_long(4278);
	dataBufferOut_long(2849) <= dataBufferIn_long(4279);
	dataBufferOut_long(3592) <= dataBufferIn_long(4280);
	dataBufferOut_long(4335) <= dataBufferIn_long(4281);
	dataBufferOut_long(5078) <= dataBufferIn_long(4282);
	dataBufferOut_long(5821) <= dataBufferIn_long(4283);
	dataBufferOut_long( 420) <= dataBufferIn_long(4284);
	dataBufferOut_long(1163) <= dataBufferIn_long(4285);
	dataBufferOut_long(1906) <= dataBufferIn_long(4286);
	dataBufferOut_long(2649) <= dataBufferIn_long(4287);
	dataBufferOut_long(3392) <= dataBufferIn_long(4288);
	dataBufferOut_long(4135) <= dataBufferIn_long(4289);
	dataBufferOut_long(4878) <= dataBufferIn_long(4290);
	dataBufferOut_long(5621) <= dataBufferIn_long(4291);
	dataBufferOut_long( 220) <= dataBufferIn_long(4292);
	dataBufferOut_long( 963) <= dataBufferIn_long(4293);
	dataBufferOut_long(1706) <= dataBufferIn_long(4294);
	dataBufferOut_long(2449) <= dataBufferIn_long(4295);
	dataBufferOut_long(3192) <= dataBufferIn_long(4296);
	dataBufferOut_long(3935) <= dataBufferIn_long(4297);
	dataBufferOut_long(4678) <= dataBufferIn_long(4298);
	dataBufferOut_long(5421) <= dataBufferIn_long(4299);
	dataBufferOut_long(  20) <= dataBufferIn_long(4300);
	dataBufferOut_long( 763) <= dataBufferIn_long(4301);
	dataBufferOut_long(1506) <= dataBufferIn_long(4302);
	dataBufferOut_long(2249) <= dataBufferIn_long(4303);
	dataBufferOut_long(2992) <= dataBufferIn_long(4304);
	dataBufferOut_long(3735) <= dataBufferIn_long(4305);
	dataBufferOut_long(4478) <= dataBufferIn_long(4306);
	dataBufferOut_long(5221) <= dataBufferIn_long(4307);
	dataBufferOut_long(5964) <= dataBufferIn_long(4308);
	dataBufferOut_long( 563) <= dataBufferIn_long(4309);
	dataBufferOut_long(1306) <= dataBufferIn_long(4310);
	dataBufferOut_long(2049) <= dataBufferIn_long(4311);
	dataBufferOut_long(2792) <= dataBufferIn_long(4312);
	dataBufferOut_long(3535) <= dataBufferIn_long(4313);
	dataBufferOut_long(4278) <= dataBufferIn_long(4314);
	dataBufferOut_long(5021) <= dataBufferIn_long(4315);
	dataBufferOut_long(5764) <= dataBufferIn_long(4316);
	dataBufferOut_long( 363) <= dataBufferIn_long(4317);
	dataBufferOut_long(1106) <= dataBufferIn_long(4318);
	dataBufferOut_long(1849) <= dataBufferIn_long(4319);
	dataBufferOut_long(2592) <= dataBufferIn_long(4320);
	dataBufferOut_long(3335) <= dataBufferIn_long(4321);
	dataBufferOut_long(4078) <= dataBufferIn_long(4322);
	dataBufferOut_long(4821) <= dataBufferIn_long(4323);
	dataBufferOut_long(5564) <= dataBufferIn_long(4324);
	dataBufferOut_long( 163) <= dataBufferIn_long(4325);
	dataBufferOut_long( 906) <= dataBufferIn_long(4326);
	dataBufferOut_long(1649) <= dataBufferIn_long(4327);
	dataBufferOut_long(2392) <= dataBufferIn_long(4328);
	dataBufferOut_long(3135) <= dataBufferIn_long(4329);
	dataBufferOut_long(3878) <= dataBufferIn_long(4330);
	dataBufferOut_long(4621) <= dataBufferIn_long(4331);
	dataBufferOut_long(5364) <= dataBufferIn_long(4332);
	dataBufferOut_long(6107) <= dataBufferIn_long(4333);
	dataBufferOut_long( 706) <= dataBufferIn_long(4334);
	dataBufferOut_long(1449) <= dataBufferIn_long(4335);
	dataBufferOut_long(2192) <= dataBufferIn_long(4336);
	dataBufferOut_long(2935) <= dataBufferIn_long(4337);
	dataBufferOut_long(3678) <= dataBufferIn_long(4338);
	dataBufferOut_long(4421) <= dataBufferIn_long(4339);
	dataBufferOut_long(5164) <= dataBufferIn_long(4340);
	dataBufferOut_long(5907) <= dataBufferIn_long(4341);
	dataBufferOut_long( 506) <= dataBufferIn_long(4342);
	dataBufferOut_long(1249) <= dataBufferIn_long(4343);
	dataBufferOut_long(1992) <= dataBufferIn_long(4344);
	dataBufferOut_long(2735) <= dataBufferIn_long(4345);
	dataBufferOut_long(3478) <= dataBufferIn_long(4346);
	dataBufferOut_long(4221) <= dataBufferIn_long(4347);
	dataBufferOut_long(4964) <= dataBufferIn_long(4348);
	dataBufferOut_long(5707) <= dataBufferIn_long(4349);
	dataBufferOut_long( 306) <= dataBufferIn_long(4350);
	dataBufferOut_long(1049) <= dataBufferIn_long(4351);
	dataBufferOut_long(1792) <= dataBufferIn_long(4352);
	dataBufferOut_long(2535) <= dataBufferIn_long(4353);
	dataBufferOut_long(3278) <= dataBufferIn_long(4354);
	dataBufferOut_long(4021) <= dataBufferIn_long(4355);
	dataBufferOut_long(4764) <= dataBufferIn_long(4356);
	dataBufferOut_long(5507) <= dataBufferIn_long(4357);
	dataBufferOut_long( 106) <= dataBufferIn_long(4358);
	dataBufferOut_long( 849) <= dataBufferIn_long(4359);
	dataBufferOut_long(1592) <= dataBufferIn_long(4360);
	dataBufferOut_long(2335) <= dataBufferIn_long(4361);
	dataBufferOut_long(3078) <= dataBufferIn_long(4362);
	dataBufferOut_long(3821) <= dataBufferIn_long(4363);
	dataBufferOut_long(4564) <= dataBufferIn_long(4364);
	dataBufferOut_long(5307) <= dataBufferIn_long(4365);
	dataBufferOut_long(6050) <= dataBufferIn_long(4366);
	dataBufferOut_long( 649) <= dataBufferIn_long(4367);
	dataBufferOut_long(1392) <= dataBufferIn_long(4368);
	dataBufferOut_long(2135) <= dataBufferIn_long(4369);
	dataBufferOut_long(2878) <= dataBufferIn_long(4370);
	dataBufferOut_long(3621) <= dataBufferIn_long(4371);
	dataBufferOut_long(4364) <= dataBufferIn_long(4372);
	dataBufferOut_long(5107) <= dataBufferIn_long(4373);
	dataBufferOut_long(5850) <= dataBufferIn_long(4374);
	dataBufferOut_long( 449) <= dataBufferIn_long(4375);
	dataBufferOut_long(1192) <= dataBufferIn_long(4376);
	dataBufferOut_long(1935) <= dataBufferIn_long(4377);
	dataBufferOut_long(2678) <= dataBufferIn_long(4378);
	dataBufferOut_long(3421) <= dataBufferIn_long(4379);
	dataBufferOut_long(4164) <= dataBufferIn_long(4380);
	dataBufferOut_long(4907) <= dataBufferIn_long(4381);
	dataBufferOut_long(5650) <= dataBufferIn_long(4382);
	dataBufferOut_long( 249) <= dataBufferIn_long(4383);
	dataBufferOut_long( 992) <= dataBufferIn_long(4384);
	dataBufferOut_long(1735) <= dataBufferIn_long(4385);
	dataBufferOut_long(2478) <= dataBufferIn_long(4386);
	dataBufferOut_long(3221) <= dataBufferIn_long(4387);
	dataBufferOut_long(3964) <= dataBufferIn_long(4388);
	dataBufferOut_long(4707) <= dataBufferIn_long(4389);
	dataBufferOut_long(5450) <= dataBufferIn_long(4390);
	dataBufferOut_long(  49) <= dataBufferIn_long(4391);
	dataBufferOut_long( 792) <= dataBufferIn_long(4392);
	dataBufferOut_long(1535) <= dataBufferIn_long(4393);
	dataBufferOut_long(2278) <= dataBufferIn_long(4394);
	dataBufferOut_long(3021) <= dataBufferIn_long(4395);
	dataBufferOut_long(3764) <= dataBufferIn_long(4396);
	dataBufferOut_long(4507) <= dataBufferIn_long(4397);
	dataBufferOut_long(5250) <= dataBufferIn_long(4398);
	dataBufferOut_long(5993) <= dataBufferIn_long(4399);
	dataBufferOut_long( 592) <= dataBufferIn_long(4400);
	dataBufferOut_long(1335) <= dataBufferIn_long(4401);
	dataBufferOut_long(2078) <= dataBufferIn_long(4402);
	dataBufferOut_long(2821) <= dataBufferIn_long(4403);
	dataBufferOut_long(3564) <= dataBufferIn_long(4404);
	dataBufferOut_long(4307) <= dataBufferIn_long(4405);
	dataBufferOut_long(5050) <= dataBufferIn_long(4406);
	dataBufferOut_long(5793) <= dataBufferIn_long(4407);
	dataBufferOut_long( 392) <= dataBufferIn_long(4408);
	dataBufferOut_long(1135) <= dataBufferIn_long(4409);
	dataBufferOut_long(1878) <= dataBufferIn_long(4410);
	dataBufferOut_long(2621) <= dataBufferIn_long(4411);
	dataBufferOut_long(3364) <= dataBufferIn_long(4412);
	dataBufferOut_long(4107) <= dataBufferIn_long(4413);
	dataBufferOut_long(4850) <= dataBufferIn_long(4414);
	dataBufferOut_long(5593) <= dataBufferIn_long(4415);
	dataBufferOut_long( 192) <= dataBufferIn_long(4416);
	dataBufferOut_long( 935) <= dataBufferIn_long(4417);
	dataBufferOut_long(1678) <= dataBufferIn_long(4418);
	dataBufferOut_long(2421) <= dataBufferIn_long(4419);
	dataBufferOut_long(3164) <= dataBufferIn_long(4420);
	dataBufferOut_long(3907) <= dataBufferIn_long(4421);
	dataBufferOut_long(4650) <= dataBufferIn_long(4422);
	dataBufferOut_long(5393) <= dataBufferIn_long(4423);
	dataBufferOut_long(6136) <= dataBufferIn_long(4424);
	dataBufferOut_long( 735) <= dataBufferIn_long(4425);
	dataBufferOut_long(1478) <= dataBufferIn_long(4426);
	dataBufferOut_long(2221) <= dataBufferIn_long(4427);
	dataBufferOut_long(2964) <= dataBufferIn_long(4428);
	dataBufferOut_long(3707) <= dataBufferIn_long(4429);
	dataBufferOut_long(4450) <= dataBufferIn_long(4430);
	dataBufferOut_long(5193) <= dataBufferIn_long(4431);
	dataBufferOut_long(5936) <= dataBufferIn_long(4432);
	dataBufferOut_long( 535) <= dataBufferIn_long(4433);
	dataBufferOut_long(1278) <= dataBufferIn_long(4434);
	dataBufferOut_long(2021) <= dataBufferIn_long(4435);
	dataBufferOut_long(2764) <= dataBufferIn_long(4436);
	dataBufferOut_long(3507) <= dataBufferIn_long(4437);
	dataBufferOut_long(4250) <= dataBufferIn_long(4438);
	dataBufferOut_long(4993) <= dataBufferIn_long(4439);
	dataBufferOut_long(5736) <= dataBufferIn_long(4440);
	dataBufferOut_long( 335) <= dataBufferIn_long(4441);
	dataBufferOut_long(1078) <= dataBufferIn_long(4442);
	dataBufferOut_long(1821) <= dataBufferIn_long(4443);
	dataBufferOut_long(2564) <= dataBufferIn_long(4444);
	dataBufferOut_long(3307) <= dataBufferIn_long(4445);
	dataBufferOut_long(4050) <= dataBufferIn_long(4446);
	dataBufferOut_long(4793) <= dataBufferIn_long(4447);
	dataBufferOut_long(5536) <= dataBufferIn_long(4448);
	dataBufferOut_long( 135) <= dataBufferIn_long(4449);
	dataBufferOut_long( 878) <= dataBufferIn_long(4450);
	dataBufferOut_long(1621) <= dataBufferIn_long(4451);
	dataBufferOut_long(2364) <= dataBufferIn_long(4452);
	dataBufferOut_long(3107) <= dataBufferIn_long(4453);
	dataBufferOut_long(3850) <= dataBufferIn_long(4454);
	dataBufferOut_long(4593) <= dataBufferIn_long(4455);
	dataBufferOut_long(5336) <= dataBufferIn_long(4456);
	dataBufferOut_long(6079) <= dataBufferIn_long(4457);
	dataBufferOut_long( 678) <= dataBufferIn_long(4458);
	dataBufferOut_long(1421) <= dataBufferIn_long(4459);
	dataBufferOut_long(2164) <= dataBufferIn_long(4460);
	dataBufferOut_long(2907) <= dataBufferIn_long(4461);
	dataBufferOut_long(3650) <= dataBufferIn_long(4462);
	dataBufferOut_long(4393) <= dataBufferIn_long(4463);
	dataBufferOut_long(5136) <= dataBufferIn_long(4464);
	dataBufferOut_long(5879) <= dataBufferIn_long(4465);
	dataBufferOut_long( 478) <= dataBufferIn_long(4466);
	dataBufferOut_long(1221) <= dataBufferIn_long(4467);
	dataBufferOut_long(1964) <= dataBufferIn_long(4468);
	dataBufferOut_long(2707) <= dataBufferIn_long(4469);
	dataBufferOut_long(3450) <= dataBufferIn_long(4470);
	dataBufferOut_long(4193) <= dataBufferIn_long(4471);
	dataBufferOut_long(4936) <= dataBufferIn_long(4472);
	dataBufferOut_long(5679) <= dataBufferIn_long(4473);
	dataBufferOut_long( 278) <= dataBufferIn_long(4474);
	dataBufferOut_long(1021) <= dataBufferIn_long(4475);
	dataBufferOut_long(1764) <= dataBufferIn_long(4476);
	dataBufferOut_long(2507) <= dataBufferIn_long(4477);
	dataBufferOut_long(3250) <= dataBufferIn_long(4478);
	dataBufferOut_long(3993) <= dataBufferIn_long(4479);
	dataBufferOut_long(4736) <= dataBufferIn_long(4480);
	dataBufferOut_long(5479) <= dataBufferIn_long(4481);
	dataBufferOut_long(  78) <= dataBufferIn_long(4482);
	dataBufferOut_long( 821) <= dataBufferIn_long(4483);
	dataBufferOut_long(1564) <= dataBufferIn_long(4484);
	dataBufferOut_long(2307) <= dataBufferIn_long(4485);
	dataBufferOut_long(3050) <= dataBufferIn_long(4486);
	dataBufferOut_long(3793) <= dataBufferIn_long(4487);
	dataBufferOut_long(4536) <= dataBufferIn_long(4488);
	dataBufferOut_long(5279) <= dataBufferIn_long(4489);
	dataBufferOut_long(6022) <= dataBufferIn_long(4490);
	dataBufferOut_long( 621) <= dataBufferIn_long(4491);
	dataBufferOut_long(1364) <= dataBufferIn_long(4492);
	dataBufferOut_long(2107) <= dataBufferIn_long(4493);
	dataBufferOut_long(2850) <= dataBufferIn_long(4494);
	dataBufferOut_long(3593) <= dataBufferIn_long(4495);
	dataBufferOut_long(4336) <= dataBufferIn_long(4496);
	dataBufferOut_long(5079) <= dataBufferIn_long(4497);
	dataBufferOut_long(5822) <= dataBufferIn_long(4498);
	dataBufferOut_long( 421) <= dataBufferIn_long(4499);
	dataBufferOut_long(1164) <= dataBufferIn_long(4500);
	dataBufferOut_long(1907) <= dataBufferIn_long(4501);
	dataBufferOut_long(2650) <= dataBufferIn_long(4502);
	dataBufferOut_long(3393) <= dataBufferIn_long(4503);
	dataBufferOut_long(4136) <= dataBufferIn_long(4504);
	dataBufferOut_long(4879) <= dataBufferIn_long(4505);
	dataBufferOut_long(5622) <= dataBufferIn_long(4506);
	dataBufferOut_long( 221) <= dataBufferIn_long(4507);
	dataBufferOut_long( 964) <= dataBufferIn_long(4508);
	dataBufferOut_long(1707) <= dataBufferIn_long(4509);
	dataBufferOut_long(2450) <= dataBufferIn_long(4510);
	dataBufferOut_long(3193) <= dataBufferIn_long(4511);
	dataBufferOut_long(3936) <= dataBufferIn_long(4512);
	dataBufferOut_long(4679) <= dataBufferIn_long(4513);
	dataBufferOut_long(5422) <= dataBufferIn_long(4514);
	dataBufferOut_long(  21) <= dataBufferIn_long(4515);
	dataBufferOut_long( 764) <= dataBufferIn_long(4516);
	dataBufferOut_long(1507) <= dataBufferIn_long(4517);
	dataBufferOut_long(2250) <= dataBufferIn_long(4518);
	dataBufferOut_long(2993) <= dataBufferIn_long(4519);
	dataBufferOut_long(3736) <= dataBufferIn_long(4520);
	dataBufferOut_long(4479) <= dataBufferIn_long(4521);
	dataBufferOut_long(5222) <= dataBufferIn_long(4522);
	dataBufferOut_long(5965) <= dataBufferIn_long(4523);
	dataBufferOut_long( 564) <= dataBufferIn_long(4524);
	dataBufferOut_long(1307) <= dataBufferIn_long(4525);
	dataBufferOut_long(2050) <= dataBufferIn_long(4526);
	dataBufferOut_long(2793) <= dataBufferIn_long(4527);
	dataBufferOut_long(3536) <= dataBufferIn_long(4528);
	dataBufferOut_long(4279) <= dataBufferIn_long(4529);
	dataBufferOut_long(5022) <= dataBufferIn_long(4530);
	dataBufferOut_long(5765) <= dataBufferIn_long(4531);
	dataBufferOut_long( 364) <= dataBufferIn_long(4532);
	dataBufferOut_long(1107) <= dataBufferIn_long(4533);
	dataBufferOut_long(1850) <= dataBufferIn_long(4534);
	dataBufferOut_long(2593) <= dataBufferIn_long(4535);
	dataBufferOut_long(3336) <= dataBufferIn_long(4536);
	dataBufferOut_long(4079) <= dataBufferIn_long(4537);
	dataBufferOut_long(4822) <= dataBufferIn_long(4538);
	dataBufferOut_long(5565) <= dataBufferIn_long(4539);
	dataBufferOut_long( 164) <= dataBufferIn_long(4540);
	dataBufferOut_long( 907) <= dataBufferIn_long(4541);
	dataBufferOut_long(1650) <= dataBufferIn_long(4542);
	dataBufferOut_long(2393) <= dataBufferIn_long(4543);
	dataBufferOut_long(3136) <= dataBufferIn_long(4544);
	dataBufferOut_long(3879) <= dataBufferIn_long(4545);
	dataBufferOut_long(4622) <= dataBufferIn_long(4546);
	dataBufferOut_long(5365) <= dataBufferIn_long(4547);
	dataBufferOut_long(6108) <= dataBufferIn_long(4548);
	dataBufferOut_long( 707) <= dataBufferIn_long(4549);
	dataBufferOut_long(1450) <= dataBufferIn_long(4550);
	dataBufferOut_long(2193) <= dataBufferIn_long(4551);
	dataBufferOut_long(2936) <= dataBufferIn_long(4552);
	dataBufferOut_long(3679) <= dataBufferIn_long(4553);
	dataBufferOut_long(4422) <= dataBufferIn_long(4554);
	dataBufferOut_long(5165) <= dataBufferIn_long(4555);
	dataBufferOut_long(5908) <= dataBufferIn_long(4556);
	dataBufferOut_long( 507) <= dataBufferIn_long(4557);
	dataBufferOut_long(1250) <= dataBufferIn_long(4558);
	dataBufferOut_long(1993) <= dataBufferIn_long(4559);
	dataBufferOut_long(2736) <= dataBufferIn_long(4560);
	dataBufferOut_long(3479) <= dataBufferIn_long(4561);
	dataBufferOut_long(4222) <= dataBufferIn_long(4562);
	dataBufferOut_long(4965) <= dataBufferIn_long(4563);
	dataBufferOut_long(5708) <= dataBufferIn_long(4564);
	dataBufferOut_long( 307) <= dataBufferIn_long(4565);
	dataBufferOut_long(1050) <= dataBufferIn_long(4566);
	dataBufferOut_long(1793) <= dataBufferIn_long(4567);
	dataBufferOut_long(2536) <= dataBufferIn_long(4568);
	dataBufferOut_long(3279) <= dataBufferIn_long(4569);
	dataBufferOut_long(4022) <= dataBufferIn_long(4570);
	dataBufferOut_long(4765) <= dataBufferIn_long(4571);
	dataBufferOut_long(5508) <= dataBufferIn_long(4572);
	dataBufferOut_long( 107) <= dataBufferIn_long(4573);
	dataBufferOut_long( 850) <= dataBufferIn_long(4574);
	dataBufferOut_long(1593) <= dataBufferIn_long(4575);
	dataBufferOut_long(2336) <= dataBufferIn_long(4576);
	dataBufferOut_long(3079) <= dataBufferIn_long(4577);
	dataBufferOut_long(3822) <= dataBufferIn_long(4578);
	dataBufferOut_long(4565) <= dataBufferIn_long(4579);
	dataBufferOut_long(5308) <= dataBufferIn_long(4580);
	dataBufferOut_long(6051) <= dataBufferIn_long(4581);
	dataBufferOut_long( 650) <= dataBufferIn_long(4582);
	dataBufferOut_long(1393) <= dataBufferIn_long(4583);
	dataBufferOut_long(2136) <= dataBufferIn_long(4584);
	dataBufferOut_long(2879) <= dataBufferIn_long(4585);
	dataBufferOut_long(3622) <= dataBufferIn_long(4586);
	dataBufferOut_long(4365) <= dataBufferIn_long(4587);
	dataBufferOut_long(5108) <= dataBufferIn_long(4588);
	dataBufferOut_long(5851) <= dataBufferIn_long(4589);
	dataBufferOut_long( 450) <= dataBufferIn_long(4590);
	dataBufferOut_long(1193) <= dataBufferIn_long(4591);
	dataBufferOut_long(1936) <= dataBufferIn_long(4592);
	dataBufferOut_long(2679) <= dataBufferIn_long(4593);
	dataBufferOut_long(3422) <= dataBufferIn_long(4594);
	dataBufferOut_long(4165) <= dataBufferIn_long(4595);
	dataBufferOut_long(4908) <= dataBufferIn_long(4596);
	dataBufferOut_long(5651) <= dataBufferIn_long(4597);
	dataBufferOut_long( 250) <= dataBufferIn_long(4598);
	dataBufferOut_long( 993) <= dataBufferIn_long(4599);
	dataBufferOut_long(1736) <= dataBufferIn_long(4600);
	dataBufferOut_long(2479) <= dataBufferIn_long(4601);
	dataBufferOut_long(3222) <= dataBufferIn_long(4602);
	dataBufferOut_long(3965) <= dataBufferIn_long(4603);
	dataBufferOut_long(4708) <= dataBufferIn_long(4604);
	dataBufferOut_long(5451) <= dataBufferIn_long(4605);
	dataBufferOut_long(  50) <= dataBufferIn_long(4606);
	dataBufferOut_long( 793) <= dataBufferIn_long(4607);
	dataBufferOut_long(1536) <= dataBufferIn_long(4608);
	dataBufferOut_long(2279) <= dataBufferIn_long(4609);
	dataBufferOut_long(3022) <= dataBufferIn_long(4610);
	dataBufferOut_long(3765) <= dataBufferIn_long(4611);
	dataBufferOut_long(4508) <= dataBufferIn_long(4612);
	dataBufferOut_long(5251) <= dataBufferIn_long(4613);
	dataBufferOut_long(5994) <= dataBufferIn_long(4614);
	dataBufferOut_long( 593) <= dataBufferIn_long(4615);
	dataBufferOut_long(1336) <= dataBufferIn_long(4616);
	dataBufferOut_long(2079) <= dataBufferIn_long(4617);
	dataBufferOut_long(2822) <= dataBufferIn_long(4618);
	dataBufferOut_long(3565) <= dataBufferIn_long(4619);
	dataBufferOut_long(4308) <= dataBufferIn_long(4620);
	dataBufferOut_long(5051) <= dataBufferIn_long(4621);
	dataBufferOut_long(5794) <= dataBufferIn_long(4622);
	dataBufferOut_long( 393) <= dataBufferIn_long(4623);
	dataBufferOut_long(1136) <= dataBufferIn_long(4624);
	dataBufferOut_long(1879) <= dataBufferIn_long(4625);
	dataBufferOut_long(2622) <= dataBufferIn_long(4626);
	dataBufferOut_long(3365) <= dataBufferIn_long(4627);
	dataBufferOut_long(4108) <= dataBufferIn_long(4628);
	dataBufferOut_long(4851) <= dataBufferIn_long(4629);
	dataBufferOut_long(5594) <= dataBufferIn_long(4630);
	dataBufferOut_long( 193) <= dataBufferIn_long(4631);
	dataBufferOut_long( 936) <= dataBufferIn_long(4632);
	dataBufferOut_long(1679) <= dataBufferIn_long(4633);
	dataBufferOut_long(2422) <= dataBufferIn_long(4634);
	dataBufferOut_long(3165) <= dataBufferIn_long(4635);
	dataBufferOut_long(3908) <= dataBufferIn_long(4636);
	dataBufferOut_long(4651) <= dataBufferIn_long(4637);
	dataBufferOut_long(5394) <= dataBufferIn_long(4638);
	dataBufferOut_long(6137) <= dataBufferIn_long(4639);
	dataBufferOut_long( 736) <= dataBufferIn_long(4640);
	dataBufferOut_long(1479) <= dataBufferIn_long(4641);
	dataBufferOut_long(2222) <= dataBufferIn_long(4642);
	dataBufferOut_long(2965) <= dataBufferIn_long(4643);
	dataBufferOut_long(3708) <= dataBufferIn_long(4644);
	dataBufferOut_long(4451) <= dataBufferIn_long(4645);
	dataBufferOut_long(5194) <= dataBufferIn_long(4646);
	dataBufferOut_long(5937) <= dataBufferIn_long(4647);
	dataBufferOut_long( 536) <= dataBufferIn_long(4648);
	dataBufferOut_long(1279) <= dataBufferIn_long(4649);
	dataBufferOut_long(2022) <= dataBufferIn_long(4650);
	dataBufferOut_long(2765) <= dataBufferIn_long(4651);
	dataBufferOut_long(3508) <= dataBufferIn_long(4652);
	dataBufferOut_long(4251) <= dataBufferIn_long(4653);
	dataBufferOut_long(4994) <= dataBufferIn_long(4654);
	dataBufferOut_long(5737) <= dataBufferIn_long(4655);
	dataBufferOut_long( 336) <= dataBufferIn_long(4656);
	dataBufferOut_long(1079) <= dataBufferIn_long(4657);
	dataBufferOut_long(1822) <= dataBufferIn_long(4658);
	dataBufferOut_long(2565) <= dataBufferIn_long(4659);
	dataBufferOut_long(3308) <= dataBufferIn_long(4660);
	dataBufferOut_long(4051) <= dataBufferIn_long(4661);
	dataBufferOut_long(4794) <= dataBufferIn_long(4662);
	dataBufferOut_long(5537) <= dataBufferIn_long(4663);
	dataBufferOut_long( 136) <= dataBufferIn_long(4664);
	dataBufferOut_long( 879) <= dataBufferIn_long(4665);
	dataBufferOut_long(1622) <= dataBufferIn_long(4666);
	dataBufferOut_long(2365) <= dataBufferIn_long(4667);
	dataBufferOut_long(3108) <= dataBufferIn_long(4668);
	dataBufferOut_long(3851) <= dataBufferIn_long(4669);
	dataBufferOut_long(4594) <= dataBufferIn_long(4670);
	dataBufferOut_long(5337) <= dataBufferIn_long(4671);
	dataBufferOut_long(6080) <= dataBufferIn_long(4672);
	dataBufferOut_long( 679) <= dataBufferIn_long(4673);
	dataBufferOut_long(1422) <= dataBufferIn_long(4674);
	dataBufferOut_long(2165) <= dataBufferIn_long(4675);
	dataBufferOut_long(2908) <= dataBufferIn_long(4676);
	dataBufferOut_long(3651) <= dataBufferIn_long(4677);
	dataBufferOut_long(4394) <= dataBufferIn_long(4678);
	dataBufferOut_long(5137) <= dataBufferIn_long(4679);
	dataBufferOut_long(5880) <= dataBufferIn_long(4680);
	dataBufferOut_long( 479) <= dataBufferIn_long(4681);
	dataBufferOut_long(1222) <= dataBufferIn_long(4682);
	dataBufferOut_long(1965) <= dataBufferIn_long(4683);
	dataBufferOut_long(2708) <= dataBufferIn_long(4684);
	dataBufferOut_long(3451) <= dataBufferIn_long(4685);
	dataBufferOut_long(4194) <= dataBufferIn_long(4686);
	dataBufferOut_long(4937) <= dataBufferIn_long(4687);
	dataBufferOut_long(5680) <= dataBufferIn_long(4688);
	dataBufferOut_long( 279) <= dataBufferIn_long(4689);
	dataBufferOut_long(1022) <= dataBufferIn_long(4690);
	dataBufferOut_long(1765) <= dataBufferIn_long(4691);
	dataBufferOut_long(2508) <= dataBufferIn_long(4692);
	dataBufferOut_long(3251) <= dataBufferIn_long(4693);
	dataBufferOut_long(3994) <= dataBufferIn_long(4694);
	dataBufferOut_long(4737) <= dataBufferIn_long(4695);
	dataBufferOut_long(5480) <= dataBufferIn_long(4696);
	dataBufferOut_long(  79) <= dataBufferIn_long(4697);
	dataBufferOut_long( 822) <= dataBufferIn_long(4698);
	dataBufferOut_long(1565) <= dataBufferIn_long(4699);
	dataBufferOut_long(2308) <= dataBufferIn_long(4700);
	dataBufferOut_long(3051) <= dataBufferIn_long(4701);
	dataBufferOut_long(3794) <= dataBufferIn_long(4702);
	dataBufferOut_long(4537) <= dataBufferIn_long(4703);
	dataBufferOut_long(5280) <= dataBufferIn_long(4704);
	dataBufferOut_long(6023) <= dataBufferIn_long(4705);
	dataBufferOut_long( 622) <= dataBufferIn_long(4706);
	dataBufferOut_long(1365) <= dataBufferIn_long(4707);
	dataBufferOut_long(2108) <= dataBufferIn_long(4708);
	dataBufferOut_long(2851) <= dataBufferIn_long(4709);
	dataBufferOut_long(3594) <= dataBufferIn_long(4710);
	dataBufferOut_long(4337) <= dataBufferIn_long(4711);
	dataBufferOut_long(5080) <= dataBufferIn_long(4712);
	dataBufferOut_long(5823) <= dataBufferIn_long(4713);
	dataBufferOut_long( 422) <= dataBufferIn_long(4714);
	dataBufferOut_long(1165) <= dataBufferIn_long(4715);
	dataBufferOut_long(1908) <= dataBufferIn_long(4716);
	dataBufferOut_long(2651) <= dataBufferIn_long(4717);
	dataBufferOut_long(3394) <= dataBufferIn_long(4718);
	dataBufferOut_long(4137) <= dataBufferIn_long(4719);
	dataBufferOut_long(4880) <= dataBufferIn_long(4720);
	dataBufferOut_long(5623) <= dataBufferIn_long(4721);
	dataBufferOut_long( 222) <= dataBufferIn_long(4722);
	dataBufferOut_long( 965) <= dataBufferIn_long(4723);
	dataBufferOut_long(1708) <= dataBufferIn_long(4724);
	dataBufferOut_long(2451) <= dataBufferIn_long(4725);
	dataBufferOut_long(3194) <= dataBufferIn_long(4726);
	dataBufferOut_long(3937) <= dataBufferIn_long(4727);
	dataBufferOut_long(4680) <= dataBufferIn_long(4728);
	dataBufferOut_long(5423) <= dataBufferIn_long(4729);
	dataBufferOut_long(  22) <= dataBufferIn_long(4730);
	dataBufferOut_long( 765) <= dataBufferIn_long(4731);
	dataBufferOut_long(1508) <= dataBufferIn_long(4732);
	dataBufferOut_long(2251) <= dataBufferIn_long(4733);
	dataBufferOut_long(2994) <= dataBufferIn_long(4734);
	dataBufferOut_long(3737) <= dataBufferIn_long(4735);
	dataBufferOut_long(4480) <= dataBufferIn_long(4736);
	dataBufferOut_long(5223) <= dataBufferIn_long(4737);
	dataBufferOut_long(5966) <= dataBufferIn_long(4738);
	dataBufferOut_long( 565) <= dataBufferIn_long(4739);
	dataBufferOut_long(1308) <= dataBufferIn_long(4740);
	dataBufferOut_long(2051) <= dataBufferIn_long(4741);
	dataBufferOut_long(2794) <= dataBufferIn_long(4742);
	dataBufferOut_long(3537) <= dataBufferIn_long(4743);
	dataBufferOut_long(4280) <= dataBufferIn_long(4744);
	dataBufferOut_long(5023) <= dataBufferIn_long(4745);
	dataBufferOut_long(5766) <= dataBufferIn_long(4746);
	dataBufferOut_long( 365) <= dataBufferIn_long(4747);
	dataBufferOut_long(1108) <= dataBufferIn_long(4748);
	dataBufferOut_long(1851) <= dataBufferIn_long(4749);
	dataBufferOut_long(2594) <= dataBufferIn_long(4750);
	dataBufferOut_long(3337) <= dataBufferIn_long(4751);
	dataBufferOut_long(4080) <= dataBufferIn_long(4752);
	dataBufferOut_long(4823) <= dataBufferIn_long(4753);
	dataBufferOut_long(5566) <= dataBufferIn_long(4754);
	dataBufferOut_long( 165) <= dataBufferIn_long(4755);
	dataBufferOut_long( 908) <= dataBufferIn_long(4756);
	dataBufferOut_long(1651) <= dataBufferIn_long(4757);
	dataBufferOut_long(2394) <= dataBufferIn_long(4758);
	dataBufferOut_long(3137) <= dataBufferIn_long(4759);
	dataBufferOut_long(3880) <= dataBufferIn_long(4760);
	dataBufferOut_long(4623) <= dataBufferIn_long(4761);
	dataBufferOut_long(5366) <= dataBufferIn_long(4762);
	dataBufferOut_long(6109) <= dataBufferIn_long(4763);
	dataBufferOut_long( 708) <= dataBufferIn_long(4764);
	dataBufferOut_long(1451) <= dataBufferIn_long(4765);
	dataBufferOut_long(2194) <= dataBufferIn_long(4766);
	dataBufferOut_long(2937) <= dataBufferIn_long(4767);
	dataBufferOut_long(3680) <= dataBufferIn_long(4768);
	dataBufferOut_long(4423) <= dataBufferIn_long(4769);
	dataBufferOut_long(5166) <= dataBufferIn_long(4770);
	dataBufferOut_long(5909) <= dataBufferIn_long(4771);
	dataBufferOut_long( 508) <= dataBufferIn_long(4772);
	dataBufferOut_long(1251) <= dataBufferIn_long(4773);
	dataBufferOut_long(1994) <= dataBufferIn_long(4774);
	dataBufferOut_long(2737) <= dataBufferIn_long(4775);
	dataBufferOut_long(3480) <= dataBufferIn_long(4776);
	dataBufferOut_long(4223) <= dataBufferIn_long(4777);
	dataBufferOut_long(4966) <= dataBufferIn_long(4778);
	dataBufferOut_long(5709) <= dataBufferIn_long(4779);
	dataBufferOut_long( 308) <= dataBufferIn_long(4780);
	dataBufferOut_long(1051) <= dataBufferIn_long(4781);
	dataBufferOut_long(1794) <= dataBufferIn_long(4782);
	dataBufferOut_long(2537) <= dataBufferIn_long(4783);
	dataBufferOut_long(3280) <= dataBufferIn_long(4784);
	dataBufferOut_long(4023) <= dataBufferIn_long(4785);
	dataBufferOut_long(4766) <= dataBufferIn_long(4786);
	dataBufferOut_long(5509) <= dataBufferIn_long(4787);
	dataBufferOut_long( 108) <= dataBufferIn_long(4788);
	dataBufferOut_long( 851) <= dataBufferIn_long(4789);
	dataBufferOut_long(1594) <= dataBufferIn_long(4790);
	dataBufferOut_long(2337) <= dataBufferIn_long(4791);
	dataBufferOut_long(3080) <= dataBufferIn_long(4792);
	dataBufferOut_long(3823) <= dataBufferIn_long(4793);
	dataBufferOut_long(4566) <= dataBufferIn_long(4794);
	dataBufferOut_long(5309) <= dataBufferIn_long(4795);
	dataBufferOut_long(6052) <= dataBufferIn_long(4796);
	dataBufferOut_long( 651) <= dataBufferIn_long(4797);
	dataBufferOut_long(1394) <= dataBufferIn_long(4798);
	dataBufferOut_long(2137) <= dataBufferIn_long(4799);
	dataBufferOut_long(2880) <= dataBufferIn_long(4800);
	dataBufferOut_long(3623) <= dataBufferIn_long(4801);
	dataBufferOut_long(4366) <= dataBufferIn_long(4802);
	dataBufferOut_long(5109) <= dataBufferIn_long(4803);
	dataBufferOut_long(5852) <= dataBufferIn_long(4804);
	dataBufferOut_long( 451) <= dataBufferIn_long(4805);
	dataBufferOut_long(1194) <= dataBufferIn_long(4806);
	dataBufferOut_long(1937) <= dataBufferIn_long(4807);
	dataBufferOut_long(2680) <= dataBufferIn_long(4808);
	dataBufferOut_long(3423) <= dataBufferIn_long(4809);
	dataBufferOut_long(4166) <= dataBufferIn_long(4810);
	dataBufferOut_long(4909) <= dataBufferIn_long(4811);
	dataBufferOut_long(5652) <= dataBufferIn_long(4812);
	dataBufferOut_long( 251) <= dataBufferIn_long(4813);
	dataBufferOut_long( 994) <= dataBufferIn_long(4814);
	dataBufferOut_long(1737) <= dataBufferIn_long(4815);
	dataBufferOut_long(2480) <= dataBufferIn_long(4816);
	dataBufferOut_long(3223) <= dataBufferIn_long(4817);
	dataBufferOut_long(3966) <= dataBufferIn_long(4818);
	dataBufferOut_long(4709) <= dataBufferIn_long(4819);
	dataBufferOut_long(5452) <= dataBufferIn_long(4820);
	dataBufferOut_long(  51) <= dataBufferIn_long(4821);
	dataBufferOut_long( 794) <= dataBufferIn_long(4822);
	dataBufferOut_long(1537) <= dataBufferIn_long(4823);
	dataBufferOut_long(2280) <= dataBufferIn_long(4824);
	dataBufferOut_long(3023) <= dataBufferIn_long(4825);
	dataBufferOut_long(3766) <= dataBufferIn_long(4826);
	dataBufferOut_long(4509) <= dataBufferIn_long(4827);
	dataBufferOut_long(5252) <= dataBufferIn_long(4828);
	dataBufferOut_long(5995) <= dataBufferIn_long(4829);
	dataBufferOut_long( 594) <= dataBufferIn_long(4830);
	dataBufferOut_long(1337) <= dataBufferIn_long(4831);
	dataBufferOut_long(2080) <= dataBufferIn_long(4832);
	dataBufferOut_long(2823) <= dataBufferIn_long(4833);
	dataBufferOut_long(3566) <= dataBufferIn_long(4834);
	dataBufferOut_long(4309) <= dataBufferIn_long(4835);
	dataBufferOut_long(5052) <= dataBufferIn_long(4836);
	dataBufferOut_long(5795) <= dataBufferIn_long(4837);
	dataBufferOut_long( 394) <= dataBufferIn_long(4838);
	dataBufferOut_long(1137) <= dataBufferIn_long(4839);
	dataBufferOut_long(1880) <= dataBufferIn_long(4840);
	dataBufferOut_long(2623) <= dataBufferIn_long(4841);
	dataBufferOut_long(3366) <= dataBufferIn_long(4842);
	dataBufferOut_long(4109) <= dataBufferIn_long(4843);
	dataBufferOut_long(4852) <= dataBufferIn_long(4844);
	dataBufferOut_long(5595) <= dataBufferIn_long(4845);
	dataBufferOut_long( 194) <= dataBufferIn_long(4846);
	dataBufferOut_long( 937) <= dataBufferIn_long(4847);
	dataBufferOut_long(1680) <= dataBufferIn_long(4848);
	dataBufferOut_long(2423) <= dataBufferIn_long(4849);
	dataBufferOut_long(3166) <= dataBufferIn_long(4850);
	dataBufferOut_long(3909) <= dataBufferIn_long(4851);
	dataBufferOut_long(4652) <= dataBufferIn_long(4852);
	dataBufferOut_long(5395) <= dataBufferIn_long(4853);
	dataBufferOut_long(6138) <= dataBufferIn_long(4854);
	dataBufferOut_long( 737) <= dataBufferIn_long(4855);
	dataBufferOut_long(1480) <= dataBufferIn_long(4856);
	dataBufferOut_long(2223) <= dataBufferIn_long(4857);
	dataBufferOut_long(2966) <= dataBufferIn_long(4858);
	dataBufferOut_long(3709) <= dataBufferIn_long(4859);
	dataBufferOut_long(4452) <= dataBufferIn_long(4860);
	dataBufferOut_long(5195) <= dataBufferIn_long(4861);
	dataBufferOut_long(5938) <= dataBufferIn_long(4862);
	dataBufferOut_long( 537) <= dataBufferIn_long(4863);
	dataBufferOut_long(1280) <= dataBufferIn_long(4864);
	dataBufferOut_long(2023) <= dataBufferIn_long(4865);
	dataBufferOut_long(2766) <= dataBufferIn_long(4866);
	dataBufferOut_long(3509) <= dataBufferIn_long(4867);
	dataBufferOut_long(4252) <= dataBufferIn_long(4868);
	dataBufferOut_long(4995) <= dataBufferIn_long(4869);
	dataBufferOut_long(5738) <= dataBufferIn_long(4870);
	dataBufferOut_long( 337) <= dataBufferIn_long(4871);
	dataBufferOut_long(1080) <= dataBufferIn_long(4872);
	dataBufferOut_long(1823) <= dataBufferIn_long(4873);
	dataBufferOut_long(2566) <= dataBufferIn_long(4874);
	dataBufferOut_long(3309) <= dataBufferIn_long(4875);
	dataBufferOut_long(4052) <= dataBufferIn_long(4876);
	dataBufferOut_long(4795) <= dataBufferIn_long(4877);
	dataBufferOut_long(5538) <= dataBufferIn_long(4878);
	dataBufferOut_long( 137) <= dataBufferIn_long(4879);
	dataBufferOut_long( 880) <= dataBufferIn_long(4880);
	dataBufferOut_long(1623) <= dataBufferIn_long(4881);
	dataBufferOut_long(2366) <= dataBufferIn_long(4882);
	dataBufferOut_long(3109) <= dataBufferIn_long(4883);
	dataBufferOut_long(3852) <= dataBufferIn_long(4884);
	dataBufferOut_long(4595) <= dataBufferIn_long(4885);
	dataBufferOut_long(5338) <= dataBufferIn_long(4886);
	dataBufferOut_long(6081) <= dataBufferIn_long(4887);
	dataBufferOut_long( 680) <= dataBufferIn_long(4888);
	dataBufferOut_long(1423) <= dataBufferIn_long(4889);
	dataBufferOut_long(2166) <= dataBufferIn_long(4890);
	dataBufferOut_long(2909) <= dataBufferIn_long(4891);
	dataBufferOut_long(3652) <= dataBufferIn_long(4892);
	dataBufferOut_long(4395) <= dataBufferIn_long(4893);
	dataBufferOut_long(5138) <= dataBufferIn_long(4894);
	dataBufferOut_long(5881) <= dataBufferIn_long(4895);
	dataBufferOut_long( 480) <= dataBufferIn_long(4896);
	dataBufferOut_long(1223) <= dataBufferIn_long(4897);
	dataBufferOut_long(1966) <= dataBufferIn_long(4898);
	dataBufferOut_long(2709) <= dataBufferIn_long(4899);
	dataBufferOut_long(3452) <= dataBufferIn_long(4900);
	dataBufferOut_long(4195) <= dataBufferIn_long(4901);
	dataBufferOut_long(4938) <= dataBufferIn_long(4902);
	dataBufferOut_long(5681) <= dataBufferIn_long(4903);
	dataBufferOut_long( 280) <= dataBufferIn_long(4904);
	dataBufferOut_long(1023) <= dataBufferIn_long(4905);
	dataBufferOut_long(1766) <= dataBufferIn_long(4906);
	dataBufferOut_long(2509) <= dataBufferIn_long(4907);
	dataBufferOut_long(3252) <= dataBufferIn_long(4908);
	dataBufferOut_long(3995) <= dataBufferIn_long(4909);
	dataBufferOut_long(4738) <= dataBufferIn_long(4910);
	dataBufferOut_long(5481) <= dataBufferIn_long(4911);
	dataBufferOut_long(  80) <= dataBufferIn_long(4912);
	dataBufferOut_long( 823) <= dataBufferIn_long(4913);
	dataBufferOut_long(1566) <= dataBufferIn_long(4914);
	dataBufferOut_long(2309) <= dataBufferIn_long(4915);
	dataBufferOut_long(3052) <= dataBufferIn_long(4916);
	dataBufferOut_long(3795) <= dataBufferIn_long(4917);
	dataBufferOut_long(4538) <= dataBufferIn_long(4918);
	dataBufferOut_long(5281) <= dataBufferIn_long(4919);
	dataBufferOut_long(6024) <= dataBufferIn_long(4920);
	dataBufferOut_long( 623) <= dataBufferIn_long(4921);
	dataBufferOut_long(1366) <= dataBufferIn_long(4922);
	dataBufferOut_long(2109) <= dataBufferIn_long(4923);
	dataBufferOut_long(2852) <= dataBufferIn_long(4924);
	dataBufferOut_long(3595) <= dataBufferIn_long(4925);
	dataBufferOut_long(4338) <= dataBufferIn_long(4926);
	dataBufferOut_long(5081) <= dataBufferIn_long(4927);
	dataBufferOut_long(5824) <= dataBufferIn_long(4928);
	dataBufferOut_long( 423) <= dataBufferIn_long(4929);
	dataBufferOut_long(1166) <= dataBufferIn_long(4930);
	dataBufferOut_long(1909) <= dataBufferIn_long(4931);
	dataBufferOut_long(2652) <= dataBufferIn_long(4932);
	dataBufferOut_long(3395) <= dataBufferIn_long(4933);
	dataBufferOut_long(4138) <= dataBufferIn_long(4934);
	dataBufferOut_long(4881) <= dataBufferIn_long(4935);
	dataBufferOut_long(5624) <= dataBufferIn_long(4936);
	dataBufferOut_long( 223) <= dataBufferIn_long(4937);
	dataBufferOut_long( 966) <= dataBufferIn_long(4938);
	dataBufferOut_long(1709) <= dataBufferIn_long(4939);
	dataBufferOut_long(2452) <= dataBufferIn_long(4940);
	dataBufferOut_long(3195) <= dataBufferIn_long(4941);
	dataBufferOut_long(3938) <= dataBufferIn_long(4942);
	dataBufferOut_long(4681) <= dataBufferIn_long(4943);
	dataBufferOut_long(5424) <= dataBufferIn_long(4944);
	dataBufferOut_long(  23) <= dataBufferIn_long(4945);
	dataBufferOut_long( 766) <= dataBufferIn_long(4946);
	dataBufferOut_long(1509) <= dataBufferIn_long(4947);
	dataBufferOut_long(2252) <= dataBufferIn_long(4948);
	dataBufferOut_long(2995) <= dataBufferIn_long(4949);
	dataBufferOut_long(3738) <= dataBufferIn_long(4950);
	dataBufferOut_long(4481) <= dataBufferIn_long(4951);
	dataBufferOut_long(5224) <= dataBufferIn_long(4952);
	dataBufferOut_long(5967) <= dataBufferIn_long(4953);
	dataBufferOut_long( 566) <= dataBufferIn_long(4954);
	dataBufferOut_long(1309) <= dataBufferIn_long(4955);
	dataBufferOut_long(2052) <= dataBufferIn_long(4956);
	dataBufferOut_long(2795) <= dataBufferIn_long(4957);
	dataBufferOut_long(3538) <= dataBufferIn_long(4958);
	dataBufferOut_long(4281) <= dataBufferIn_long(4959);
	dataBufferOut_long(5024) <= dataBufferIn_long(4960);
	dataBufferOut_long(5767) <= dataBufferIn_long(4961);
	dataBufferOut_long( 366) <= dataBufferIn_long(4962);
	dataBufferOut_long(1109) <= dataBufferIn_long(4963);
	dataBufferOut_long(1852) <= dataBufferIn_long(4964);
	dataBufferOut_long(2595) <= dataBufferIn_long(4965);
	dataBufferOut_long(3338) <= dataBufferIn_long(4966);
	dataBufferOut_long(4081) <= dataBufferIn_long(4967);
	dataBufferOut_long(4824) <= dataBufferIn_long(4968);
	dataBufferOut_long(5567) <= dataBufferIn_long(4969);
	dataBufferOut_long( 166) <= dataBufferIn_long(4970);
	dataBufferOut_long( 909) <= dataBufferIn_long(4971);
	dataBufferOut_long(1652) <= dataBufferIn_long(4972);
	dataBufferOut_long(2395) <= dataBufferIn_long(4973);
	dataBufferOut_long(3138) <= dataBufferIn_long(4974);
	dataBufferOut_long(3881) <= dataBufferIn_long(4975);
	dataBufferOut_long(4624) <= dataBufferIn_long(4976);
	dataBufferOut_long(5367) <= dataBufferIn_long(4977);
	dataBufferOut_long(6110) <= dataBufferIn_long(4978);
	dataBufferOut_long( 709) <= dataBufferIn_long(4979);
	dataBufferOut_long(1452) <= dataBufferIn_long(4980);
	dataBufferOut_long(2195) <= dataBufferIn_long(4981);
	dataBufferOut_long(2938) <= dataBufferIn_long(4982);
	dataBufferOut_long(3681) <= dataBufferIn_long(4983);
	dataBufferOut_long(4424) <= dataBufferIn_long(4984);
	dataBufferOut_long(5167) <= dataBufferIn_long(4985);
	dataBufferOut_long(5910) <= dataBufferIn_long(4986);
	dataBufferOut_long( 509) <= dataBufferIn_long(4987);
	dataBufferOut_long(1252) <= dataBufferIn_long(4988);
	dataBufferOut_long(1995) <= dataBufferIn_long(4989);
	dataBufferOut_long(2738) <= dataBufferIn_long(4990);
	dataBufferOut_long(3481) <= dataBufferIn_long(4991);
	dataBufferOut_long(4224) <= dataBufferIn_long(4992);
	dataBufferOut_long(4967) <= dataBufferIn_long(4993);
	dataBufferOut_long(5710) <= dataBufferIn_long(4994);
	dataBufferOut_long( 309) <= dataBufferIn_long(4995);
	dataBufferOut_long(1052) <= dataBufferIn_long(4996);
	dataBufferOut_long(1795) <= dataBufferIn_long(4997);
	dataBufferOut_long(2538) <= dataBufferIn_long(4998);
	dataBufferOut_long(3281) <= dataBufferIn_long(4999);
	dataBufferOut_long(4024) <= dataBufferIn_long(5000);
	dataBufferOut_long(4767) <= dataBufferIn_long(5001);
	dataBufferOut_long(5510) <= dataBufferIn_long(5002);
	dataBufferOut_long( 109) <= dataBufferIn_long(5003);
	dataBufferOut_long( 852) <= dataBufferIn_long(5004);
	dataBufferOut_long(1595) <= dataBufferIn_long(5005);
	dataBufferOut_long(2338) <= dataBufferIn_long(5006);
	dataBufferOut_long(3081) <= dataBufferIn_long(5007);
	dataBufferOut_long(3824) <= dataBufferIn_long(5008);
	dataBufferOut_long(4567) <= dataBufferIn_long(5009);
	dataBufferOut_long(5310) <= dataBufferIn_long(5010);
	dataBufferOut_long(6053) <= dataBufferIn_long(5011);
	dataBufferOut_long( 652) <= dataBufferIn_long(5012);
	dataBufferOut_long(1395) <= dataBufferIn_long(5013);
	dataBufferOut_long(2138) <= dataBufferIn_long(5014);
	dataBufferOut_long(2881) <= dataBufferIn_long(5015);
	dataBufferOut_long(3624) <= dataBufferIn_long(5016);
	dataBufferOut_long(4367) <= dataBufferIn_long(5017);
	dataBufferOut_long(5110) <= dataBufferIn_long(5018);
	dataBufferOut_long(5853) <= dataBufferIn_long(5019);
	dataBufferOut_long( 452) <= dataBufferIn_long(5020);
	dataBufferOut_long(1195) <= dataBufferIn_long(5021);
	dataBufferOut_long(1938) <= dataBufferIn_long(5022);
	dataBufferOut_long(2681) <= dataBufferIn_long(5023);
	dataBufferOut_long(3424) <= dataBufferIn_long(5024);
	dataBufferOut_long(4167) <= dataBufferIn_long(5025);
	dataBufferOut_long(4910) <= dataBufferIn_long(5026);
	dataBufferOut_long(5653) <= dataBufferIn_long(5027);
	dataBufferOut_long( 252) <= dataBufferIn_long(5028);
	dataBufferOut_long( 995) <= dataBufferIn_long(5029);
	dataBufferOut_long(1738) <= dataBufferIn_long(5030);
	dataBufferOut_long(2481) <= dataBufferIn_long(5031);
	dataBufferOut_long(3224) <= dataBufferIn_long(5032);
	dataBufferOut_long(3967) <= dataBufferIn_long(5033);
	dataBufferOut_long(4710) <= dataBufferIn_long(5034);
	dataBufferOut_long(5453) <= dataBufferIn_long(5035);
	dataBufferOut_long(  52) <= dataBufferIn_long(5036);
	dataBufferOut_long( 795) <= dataBufferIn_long(5037);
	dataBufferOut_long(1538) <= dataBufferIn_long(5038);
	dataBufferOut_long(2281) <= dataBufferIn_long(5039);
	dataBufferOut_long(3024) <= dataBufferIn_long(5040);
	dataBufferOut_long(3767) <= dataBufferIn_long(5041);
	dataBufferOut_long(4510) <= dataBufferIn_long(5042);
	dataBufferOut_long(5253) <= dataBufferIn_long(5043);
	dataBufferOut_long(5996) <= dataBufferIn_long(5044);
	dataBufferOut_long( 595) <= dataBufferIn_long(5045);
	dataBufferOut_long(1338) <= dataBufferIn_long(5046);
	dataBufferOut_long(2081) <= dataBufferIn_long(5047);
	dataBufferOut_long(2824) <= dataBufferIn_long(5048);
	dataBufferOut_long(3567) <= dataBufferIn_long(5049);
	dataBufferOut_long(4310) <= dataBufferIn_long(5050);
	dataBufferOut_long(5053) <= dataBufferIn_long(5051);
	dataBufferOut_long(5796) <= dataBufferIn_long(5052);
	dataBufferOut_long( 395) <= dataBufferIn_long(5053);
	dataBufferOut_long(1138) <= dataBufferIn_long(5054);
	dataBufferOut_long(1881) <= dataBufferIn_long(5055);
	dataBufferOut_long(2624) <= dataBufferIn_long(5056);
	dataBufferOut_long(3367) <= dataBufferIn_long(5057);
	dataBufferOut_long(4110) <= dataBufferIn_long(5058);
	dataBufferOut_long(4853) <= dataBufferIn_long(5059);
	dataBufferOut_long(5596) <= dataBufferIn_long(5060);
	dataBufferOut_long( 195) <= dataBufferIn_long(5061);
	dataBufferOut_long( 938) <= dataBufferIn_long(5062);
	dataBufferOut_long(1681) <= dataBufferIn_long(5063);
	dataBufferOut_long(2424) <= dataBufferIn_long(5064);
	dataBufferOut_long(3167) <= dataBufferIn_long(5065);
	dataBufferOut_long(3910) <= dataBufferIn_long(5066);
	dataBufferOut_long(4653) <= dataBufferIn_long(5067);
	dataBufferOut_long(5396) <= dataBufferIn_long(5068);
	dataBufferOut_long(6139) <= dataBufferIn_long(5069);
	dataBufferOut_long( 738) <= dataBufferIn_long(5070);
	dataBufferOut_long(1481) <= dataBufferIn_long(5071);
	dataBufferOut_long(2224) <= dataBufferIn_long(5072);
	dataBufferOut_long(2967) <= dataBufferIn_long(5073);
	dataBufferOut_long(3710) <= dataBufferIn_long(5074);
	dataBufferOut_long(4453) <= dataBufferIn_long(5075);
	dataBufferOut_long(5196) <= dataBufferIn_long(5076);
	dataBufferOut_long(5939) <= dataBufferIn_long(5077);
	dataBufferOut_long( 538) <= dataBufferIn_long(5078);
	dataBufferOut_long(1281) <= dataBufferIn_long(5079);
	dataBufferOut_long(2024) <= dataBufferIn_long(5080);
	dataBufferOut_long(2767) <= dataBufferIn_long(5081);
	dataBufferOut_long(3510) <= dataBufferIn_long(5082);
	dataBufferOut_long(4253) <= dataBufferIn_long(5083);
	dataBufferOut_long(4996) <= dataBufferIn_long(5084);
	dataBufferOut_long(5739) <= dataBufferIn_long(5085);
	dataBufferOut_long( 338) <= dataBufferIn_long(5086);
	dataBufferOut_long(1081) <= dataBufferIn_long(5087);
	dataBufferOut_long(1824) <= dataBufferIn_long(5088);
	dataBufferOut_long(2567) <= dataBufferIn_long(5089);
	dataBufferOut_long(3310) <= dataBufferIn_long(5090);
	dataBufferOut_long(4053) <= dataBufferIn_long(5091);
	dataBufferOut_long(4796) <= dataBufferIn_long(5092);
	dataBufferOut_long(5539) <= dataBufferIn_long(5093);
	dataBufferOut_long( 138) <= dataBufferIn_long(5094);
	dataBufferOut_long( 881) <= dataBufferIn_long(5095);
	dataBufferOut_long(1624) <= dataBufferIn_long(5096);
	dataBufferOut_long(2367) <= dataBufferIn_long(5097);
	dataBufferOut_long(3110) <= dataBufferIn_long(5098);
	dataBufferOut_long(3853) <= dataBufferIn_long(5099);
	dataBufferOut_long(4596) <= dataBufferIn_long(5100);
	dataBufferOut_long(5339) <= dataBufferIn_long(5101);
	dataBufferOut_long(6082) <= dataBufferIn_long(5102);
	dataBufferOut_long( 681) <= dataBufferIn_long(5103);
	dataBufferOut_long(1424) <= dataBufferIn_long(5104);
	dataBufferOut_long(2167) <= dataBufferIn_long(5105);
	dataBufferOut_long(2910) <= dataBufferIn_long(5106);
	dataBufferOut_long(3653) <= dataBufferIn_long(5107);
	dataBufferOut_long(4396) <= dataBufferIn_long(5108);
	dataBufferOut_long(5139) <= dataBufferIn_long(5109);
	dataBufferOut_long(5882) <= dataBufferIn_long(5110);
	dataBufferOut_long( 481) <= dataBufferIn_long(5111);
	dataBufferOut_long(1224) <= dataBufferIn_long(5112);
	dataBufferOut_long(1967) <= dataBufferIn_long(5113);
	dataBufferOut_long(2710) <= dataBufferIn_long(5114);
	dataBufferOut_long(3453) <= dataBufferIn_long(5115);
	dataBufferOut_long(4196) <= dataBufferIn_long(5116);
	dataBufferOut_long(4939) <= dataBufferIn_long(5117);
	dataBufferOut_long(5682) <= dataBufferIn_long(5118);
	dataBufferOut_long( 281) <= dataBufferIn_long(5119);
	dataBufferOut_long(1024) <= dataBufferIn_long(5120);
	dataBufferOut_long(1767) <= dataBufferIn_long(5121);
	dataBufferOut_long(2510) <= dataBufferIn_long(5122);
	dataBufferOut_long(3253) <= dataBufferIn_long(5123);
	dataBufferOut_long(3996) <= dataBufferIn_long(5124);
	dataBufferOut_long(4739) <= dataBufferIn_long(5125);
	dataBufferOut_long(5482) <= dataBufferIn_long(5126);
	dataBufferOut_long(  81) <= dataBufferIn_long(5127);
	dataBufferOut_long( 824) <= dataBufferIn_long(5128);
	dataBufferOut_long(1567) <= dataBufferIn_long(5129);
	dataBufferOut_long(2310) <= dataBufferIn_long(5130);
	dataBufferOut_long(3053) <= dataBufferIn_long(5131);
	dataBufferOut_long(3796) <= dataBufferIn_long(5132);
	dataBufferOut_long(4539) <= dataBufferIn_long(5133);
	dataBufferOut_long(5282) <= dataBufferIn_long(5134);
	dataBufferOut_long(6025) <= dataBufferIn_long(5135);
	dataBufferOut_long( 624) <= dataBufferIn_long(5136);
	dataBufferOut_long(1367) <= dataBufferIn_long(5137);
	dataBufferOut_long(2110) <= dataBufferIn_long(5138);
	dataBufferOut_long(2853) <= dataBufferIn_long(5139);
	dataBufferOut_long(3596) <= dataBufferIn_long(5140);
	dataBufferOut_long(4339) <= dataBufferIn_long(5141);
	dataBufferOut_long(5082) <= dataBufferIn_long(5142);
	dataBufferOut_long(5825) <= dataBufferIn_long(5143);
	dataBufferOut_long( 424) <= dataBufferIn_long(5144);
	dataBufferOut_long(1167) <= dataBufferIn_long(5145);
	dataBufferOut_long(1910) <= dataBufferIn_long(5146);
	dataBufferOut_long(2653) <= dataBufferIn_long(5147);
	dataBufferOut_long(3396) <= dataBufferIn_long(5148);
	dataBufferOut_long(4139) <= dataBufferIn_long(5149);
	dataBufferOut_long(4882) <= dataBufferIn_long(5150);
	dataBufferOut_long(5625) <= dataBufferIn_long(5151);
	dataBufferOut_long( 224) <= dataBufferIn_long(5152);
	dataBufferOut_long( 967) <= dataBufferIn_long(5153);
	dataBufferOut_long(1710) <= dataBufferIn_long(5154);
	dataBufferOut_long(2453) <= dataBufferIn_long(5155);
	dataBufferOut_long(3196) <= dataBufferIn_long(5156);
	dataBufferOut_long(3939) <= dataBufferIn_long(5157);
	dataBufferOut_long(4682) <= dataBufferIn_long(5158);
	dataBufferOut_long(5425) <= dataBufferIn_long(5159);
	dataBufferOut_long(  24) <= dataBufferIn_long(5160);
	dataBufferOut_long( 767) <= dataBufferIn_long(5161);
	dataBufferOut_long(1510) <= dataBufferIn_long(5162);
	dataBufferOut_long(2253) <= dataBufferIn_long(5163);
	dataBufferOut_long(2996) <= dataBufferIn_long(5164);
	dataBufferOut_long(3739) <= dataBufferIn_long(5165);
	dataBufferOut_long(4482) <= dataBufferIn_long(5166);
	dataBufferOut_long(5225) <= dataBufferIn_long(5167);
	dataBufferOut_long(5968) <= dataBufferIn_long(5168);
	dataBufferOut_long( 567) <= dataBufferIn_long(5169);
	dataBufferOut_long(1310) <= dataBufferIn_long(5170);
	dataBufferOut_long(2053) <= dataBufferIn_long(5171);
	dataBufferOut_long(2796) <= dataBufferIn_long(5172);
	dataBufferOut_long(3539) <= dataBufferIn_long(5173);
	dataBufferOut_long(4282) <= dataBufferIn_long(5174);
	dataBufferOut_long(5025) <= dataBufferIn_long(5175);
	dataBufferOut_long(5768) <= dataBufferIn_long(5176);
	dataBufferOut_long( 367) <= dataBufferIn_long(5177);
	dataBufferOut_long(1110) <= dataBufferIn_long(5178);
	dataBufferOut_long(1853) <= dataBufferIn_long(5179);
	dataBufferOut_long(2596) <= dataBufferIn_long(5180);
	dataBufferOut_long(3339) <= dataBufferIn_long(5181);
	dataBufferOut_long(4082) <= dataBufferIn_long(5182);
	dataBufferOut_long(4825) <= dataBufferIn_long(5183);
	dataBufferOut_long(5568) <= dataBufferIn_long(5184);
	dataBufferOut_long( 167) <= dataBufferIn_long(5185);
	dataBufferOut_long( 910) <= dataBufferIn_long(5186);
	dataBufferOut_long(1653) <= dataBufferIn_long(5187);
	dataBufferOut_long(2396) <= dataBufferIn_long(5188);
	dataBufferOut_long(3139) <= dataBufferIn_long(5189);
	dataBufferOut_long(3882) <= dataBufferIn_long(5190);
	dataBufferOut_long(4625) <= dataBufferIn_long(5191);
	dataBufferOut_long(5368) <= dataBufferIn_long(5192);
	dataBufferOut_long(6111) <= dataBufferIn_long(5193);
	dataBufferOut_long( 710) <= dataBufferIn_long(5194);
	dataBufferOut_long(1453) <= dataBufferIn_long(5195);
	dataBufferOut_long(2196) <= dataBufferIn_long(5196);
	dataBufferOut_long(2939) <= dataBufferIn_long(5197);
	dataBufferOut_long(3682) <= dataBufferIn_long(5198);
	dataBufferOut_long(4425) <= dataBufferIn_long(5199);
	dataBufferOut_long(5168) <= dataBufferIn_long(5200);
	dataBufferOut_long(5911) <= dataBufferIn_long(5201);
	dataBufferOut_long( 510) <= dataBufferIn_long(5202);
	dataBufferOut_long(1253) <= dataBufferIn_long(5203);
	dataBufferOut_long(1996) <= dataBufferIn_long(5204);
	dataBufferOut_long(2739) <= dataBufferIn_long(5205);
	dataBufferOut_long(3482) <= dataBufferIn_long(5206);
	dataBufferOut_long(4225) <= dataBufferIn_long(5207);
	dataBufferOut_long(4968) <= dataBufferIn_long(5208);
	dataBufferOut_long(5711) <= dataBufferIn_long(5209);
	dataBufferOut_long( 310) <= dataBufferIn_long(5210);
	dataBufferOut_long(1053) <= dataBufferIn_long(5211);
	dataBufferOut_long(1796) <= dataBufferIn_long(5212);
	dataBufferOut_long(2539) <= dataBufferIn_long(5213);
	dataBufferOut_long(3282) <= dataBufferIn_long(5214);
	dataBufferOut_long(4025) <= dataBufferIn_long(5215);
	dataBufferOut_long(4768) <= dataBufferIn_long(5216);
	dataBufferOut_long(5511) <= dataBufferIn_long(5217);
	dataBufferOut_long( 110) <= dataBufferIn_long(5218);
	dataBufferOut_long( 853) <= dataBufferIn_long(5219);
	dataBufferOut_long(1596) <= dataBufferIn_long(5220);
	dataBufferOut_long(2339) <= dataBufferIn_long(5221);
	dataBufferOut_long(3082) <= dataBufferIn_long(5222);
	dataBufferOut_long(3825) <= dataBufferIn_long(5223);
	dataBufferOut_long(4568) <= dataBufferIn_long(5224);
	dataBufferOut_long(5311) <= dataBufferIn_long(5225);
	dataBufferOut_long(6054) <= dataBufferIn_long(5226);
	dataBufferOut_long( 653) <= dataBufferIn_long(5227);
	dataBufferOut_long(1396) <= dataBufferIn_long(5228);
	dataBufferOut_long(2139) <= dataBufferIn_long(5229);
	dataBufferOut_long(2882) <= dataBufferIn_long(5230);
	dataBufferOut_long(3625) <= dataBufferIn_long(5231);
	dataBufferOut_long(4368) <= dataBufferIn_long(5232);
	dataBufferOut_long(5111) <= dataBufferIn_long(5233);
	dataBufferOut_long(5854) <= dataBufferIn_long(5234);
	dataBufferOut_long( 453) <= dataBufferIn_long(5235);
	dataBufferOut_long(1196) <= dataBufferIn_long(5236);
	dataBufferOut_long(1939) <= dataBufferIn_long(5237);
	dataBufferOut_long(2682) <= dataBufferIn_long(5238);
	dataBufferOut_long(3425) <= dataBufferIn_long(5239);
	dataBufferOut_long(4168) <= dataBufferIn_long(5240);
	dataBufferOut_long(4911) <= dataBufferIn_long(5241);
	dataBufferOut_long(5654) <= dataBufferIn_long(5242);
	dataBufferOut_long( 253) <= dataBufferIn_long(5243);
	dataBufferOut_long( 996) <= dataBufferIn_long(5244);
	dataBufferOut_long(1739) <= dataBufferIn_long(5245);
	dataBufferOut_long(2482) <= dataBufferIn_long(5246);
	dataBufferOut_long(3225) <= dataBufferIn_long(5247);
	dataBufferOut_long(3968) <= dataBufferIn_long(5248);
	dataBufferOut_long(4711) <= dataBufferIn_long(5249);
	dataBufferOut_long(5454) <= dataBufferIn_long(5250);
	dataBufferOut_long(  53) <= dataBufferIn_long(5251);
	dataBufferOut_long( 796) <= dataBufferIn_long(5252);
	dataBufferOut_long(1539) <= dataBufferIn_long(5253);
	dataBufferOut_long(2282) <= dataBufferIn_long(5254);
	dataBufferOut_long(3025) <= dataBufferIn_long(5255);
	dataBufferOut_long(3768) <= dataBufferIn_long(5256);
	dataBufferOut_long(4511) <= dataBufferIn_long(5257);
	dataBufferOut_long(5254) <= dataBufferIn_long(5258);
	dataBufferOut_long(5997) <= dataBufferIn_long(5259);
	dataBufferOut_long( 596) <= dataBufferIn_long(5260);
	dataBufferOut_long(1339) <= dataBufferIn_long(5261);
	dataBufferOut_long(2082) <= dataBufferIn_long(5262);
	dataBufferOut_long(2825) <= dataBufferIn_long(5263);
	dataBufferOut_long(3568) <= dataBufferIn_long(5264);
	dataBufferOut_long(4311) <= dataBufferIn_long(5265);
	dataBufferOut_long(5054) <= dataBufferIn_long(5266);
	dataBufferOut_long(5797) <= dataBufferIn_long(5267);
	dataBufferOut_long( 396) <= dataBufferIn_long(5268);
	dataBufferOut_long(1139) <= dataBufferIn_long(5269);
	dataBufferOut_long(1882) <= dataBufferIn_long(5270);
	dataBufferOut_long(2625) <= dataBufferIn_long(5271);
	dataBufferOut_long(3368) <= dataBufferIn_long(5272);
	dataBufferOut_long(4111) <= dataBufferIn_long(5273);
	dataBufferOut_long(4854) <= dataBufferIn_long(5274);
	dataBufferOut_long(5597) <= dataBufferIn_long(5275);
	dataBufferOut_long( 196) <= dataBufferIn_long(5276);
	dataBufferOut_long( 939) <= dataBufferIn_long(5277);
	dataBufferOut_long(1682) <= dataBufferIn_long(5278);
	dataBufferOut_long(2425) <= dataBufferIn_long(5279);
	dataBufferOut_long(3168) <= dataBufferIn_long(5280);
	dataBufferOut_long(3911) <= dataBufferIn_long(5281);
	dataBufferOut_long(4654) <= dataBufferIn_long(5282);
	dataBufferOut_long(5397) <= dataBufferIn_long(5283);
	dataBufferOut_long(6140) <= dataBufferIn_long(5284);
	dataBufferOut_long( 739) <= dataBufferIn_long(5285);
	dataBufferOut_long(1482) <= dataBufferIn_long(5286);
	dataBufferOut_long(2225) <= dataBufferIn_long(5287);
	dataBufferOut_long(2968) <= dataBufferIn_long(5288);
	dataBufferOut_long(3711) <= dataBufferIn_long(5289);
	dataBufferOut_long(4454) <= dataBufferIn_long(5290);
	dataBufferOut_long(5197) <= dataBufferIn_long(5291);
	dataBufferOut_long(5940) <= dataBufferIn_long(5292);
	dataBufferOut_long( 539) <= dataBufferIn_long(5293);
	dataBufferOut_long(1282) <= dataBufferIn_long(5294);
	dataBufferOut_long(2025) <= dataBufferIn_long(5295);
	dataBufferOut_long(2768) <= dataBufferIn_long(5296);
	dataBufferOut_long(3511) <= dataBufferIn_long(5297);
	dataBufferOut_long(4254) <= dataBufferIn_long(5298);
	dataBufferOut_long(4997) <= dataBufferIn_long(5299);
	dataBufferOut_long(5740) <= dataBufferIn_long(5300);
	dataBufferOut_long( 339) <= dataBufferIn_long(5301);
	dataBufferOut_long(1082) <= dataBufferIn_long(5302);
	dataBufferOut_long(1825) <= dataBufferIn_long(5303);
	dataBufferOut_long(2568) <= dataBufferIn_long(5304);
	dataBufferOut_long(3311) <= dataBufferIn_long(5305);
	dataBufferOut_long(4054) <= dataBufferIn_long(5306);
	dataBufferOut_long(4797) <= dataBufferIn_long(5307);
	dataBufferOut_long(5540) <= dataBufferIn_long(5308);
	dataBufferOut_long( 139) <= dataBufferIn_long(5309);
	dataBufferOut_long( 882) <= dataBufferIn_long(5310);
	dataBufferOut_long(1625) <= dataBufferIn_long(5311);
	dataBufferOut_long(2368) <= dataBufferIn_long(5312);
	dataBufferOut_long(3111) <= dataBufferIn_long(5313);
	dataBufferOut_long(3854) <= dataBufferIn_long(5314);
	dataBufferOut_long(4597) <= dataBufferIn_long(5315);
	dataBufferOut_long(5340) <= dataBufferIn_long(5316);
	dataBufferOut_long(6083) <= dataBufferIn_long(5317);
	dataBufferOut_long( 682) <= dataBufferIn_long(5318);
	dataBufferOut_long(1425) <= dataBufferIn_long(5319);
	dataBufferOut_long(2168) <= dataBufferIn_long(5320);
	dataBufferOut_long(2911) <= dataBufferIn_long(5321);
	dataBufferOut_long(3654) <= dataBufferIn_long(5322);
	dataBufferOut_long(4397) <= dataBufferIn_long(5323);
	dataBufferOut_long(5140) <= dataBufferIn_long(5324);
	dataBufferOut_long(5883) <= dataBufferIn_long(5325);
	dataBufferOut_long( 482) <= dataBufferIn_long(5326);
	dataBufferOut_long(1225) <= dataBufferIn_long(5327);
	dataBufferOut_long(1968) <= dataBufferIn_long(5328);
	dataBufferOut_long(2711) <= dataBufferIn_long(5329);
	dataBufferOut_long(3454) <= dataBufferIn_long(5330);
	dataBufferOut_long(4197) <= dataBufferIn_long(5331);
	dataBufferOut_long(4940) <= dataBufferIn_long(5332);
	dataBufferOut_long(5683) <= dataBufferIn_long(5333);
	dataBufferOut_long( 282) <= dataBufferIn_long(5334);
	dataBufferOut_long(1025) <= dataBufferIn_long(5335);
	dataBufferOut_long(1768) <= dataBufferIn_long(5336);
	dataBufferOut_long(2511) <= dataBufferIn_long(5337);
	dataBufferOut_long(3254) <= dataBufferIn_long(5338);
	dataBufferOut_long(3997) <= dataBufferIn_long(5339);
	dataBufferOut_long(4740) <= dataBufferIn_long(5340);
	dataBufferOut_long(5483) <= dataBufferIn_long(5341);
	dataBufferOut_long(  82) <= dataBufferIn_long(5342);
	dataBufferOut_long( 825) <= dataBufferIn_long(5343);
	dataBufferOut_long(1568) <= dataBufferIn_long(5344);
	dataBufferOut_long(2311) <= dataBufferIn_long(5345);
	dataBufferOut_long(3054) <= dataBufferIn_long(5346);
	dataBufferOut_long(3797) <= dataBufferIn_long(5347);
	dataBufferOut_long(4540) <= dataBufferIn_long(5348);
	dataBufferOut_long(5283) <= dataBufferIn_long(5349);
	dataBufferOut_long(6026) <= dataBufferIn_long(5350);
	dataBufferOut_long( 625) <= dataBufferIn_long(5351);
	dataBufferOut_long(1368) <= dataBufferIn_long(5352);
	dataBufferOut_long(2111) <= dataBufferIn_long(5353);
	dataBufferOut_long(2854) <= dataBufferIn_long(5354);
	dataBufferOut_long(3597) <= dataBufferIn_long(5355);
	dataBufferOut_long(4340) <= dataBufferIn_long(5356);
	dataBufferOut_long(5083) <= dataBufferIn_long(5357);
	dataBufferOut_long(5826) <= dataBufferIn_long(5358);
	dataBufferOut_long( 425) <= dataBufferIn_long(5359);
	dataBufferOut_long(1168) <= dataBufferIn_long(5360);
	dataBufferOut_long(1911) <= dataBufferIn_long(5361);
	dataBufferOut_long(2654) <= dataBufferIn_long(5362);
	dataBufferOut_long(3397) <= dataBufferIn_long(5363);
	dataBufferOut_long(4140) <= dataBufferIn_long(5364);
	dataBufferOut_long(4883) <= dataBufferIn_long(5365);
	dataBufferOut_long(5626) <= dataBufferIn_long(5366);
	dataBufferOut_long( 225) <= dataBufferIn_long(5367);
	dataBufferOut_long( 968) <= dataBufferIn_long(5368);
	dataBufferOut_long(1711) <= dataBufferIn_long(5369);
	dataBufferOut_long(2454) <= dataBufferIn_long(5370);
	dataBufferOut_long(3197) <= dataBufferIn_long(5371);
	dataBufferOut_long(3940) <= dataBufferIn_long(5372);
	dataBufferOut_long(4683) <= dataBufferIn_long(5373);
	dataBufferOut_long(5426) <= dataBufferIn_long(5374);
	dataBufferOut_long(  25) <= dataBufferIn_long(5375);
	dataBufferOut_long( 768) <= dataBufferIn_long(5376);
	dataBufferOut_long(1511) <= dataBufferIn_long(5377);
	dataBufferOut_long(2254) <= dataBufferIn_long(5378);
	dataBufferOut_long(2997) <= dataBufferIn_long(5379);
	dataBufferOut_long(3740) <= dataBufferIn_long(5380);
	dataBufferOut_long(4483) <= dataBufferIn_long(5381);
	dataBufferOut_long(5226) <= dataBufferIn_long(5382);
	dataBufferOut_long(5969) <= dataBufferIn_long(5383);
	dataBufferOut_long( 568) <= dataBufferIn_long(5384);
	dataBufferOut_long(1311) <= dataBufferIn_long(5385);
	dataBufferOut_long(2054) <= dataBufferIn_long(5386);
	dataBufferOut_long(2797) <= dataBufferIn_long(5387);
	dataBufferOut_long(3540) <= dataBufferIn_long(5388);
	dataBufferOut_long(4283) <= dataBufferIn_long(5389);
	dataBufferOut_long(5026) <= dataBufferIn_long(5390);
	dataBufferOut_long(5769) <= dataBufferIn_long(5391);
	dataBufferOut_long( 368) <= dataBufferIn_long(5392);
	dataBufferOut_long(1111) <= dataBufferIn_long(5393);
	dataBufferOut_long(1854) <= dataBufferIn_long(5394);
	dataBufferOut_long(2597) <= dataBufferIn_long(5395);
	dataBufferOut_long(3340) <= dataBufferIn_long(5396);
	dataBufferOut_long(4083) <= dataBufferIn_long(5397);
	dataBufferOut_long(4826) <= dataBufferIn_long(5398);
	dataBufferOut_long(5569) <= dataBufferIn_long(5399);
	dataBufferOut_long( 168) <= dataBufferIn_long(5400);
	dataBufferOut_long( 911) <= dataBufferIn_long(5401);
	dataBufferOut_long(1654) <= dataBufferIn_long(5402);
	dataBufferOut_long(2397) <= dataBufferIn_long(5403);
	dataBufferOut_long(3140) <= dataBufferIn_long(5404);
	dataBufferOut_long(3883) <= dataBufferIn_long(5405);
	dataBufferOut_long(4626) <= dataBufferIn_long(5406);
	dataBufferOut_long(5369) <= dataBufferIn_long(5407);
	dataBufferOut_long(6112) <= dataBufferIn_long(5408);
	dataBufferOut_long( 711) <= dataBufferIn_long(5409);
	dataBufferOut_long(1454) <= dataBufferIn_long(5410);
	dataBufferOut_long(2197) <= dataBufferIn_long(5411);
	dataBufferOut_long(2940) <= dataBufferIn_long(5412);
	dataBufferOut_long(3683) <= dataBufferIn_long(5413);
	dataBufferOut_long(4426) <= dataBufferIn_long(5414);
	dataBufferOut_long(5169) <= dataBufferIn_long(5415);
	dataBufferOut_long(5912) <= dataBufferIn_long(5416);
	dataBufferOut_long( 511) <= dataBufferIn_long(5417);
	dataBufferOut_long(1254) <= dataBufferIn_long(5418);
	dataBufferOut_long(1997) <= dataBufferIn_long(5419);
	dataBufferOut_long(2740) <= dataBufferIn_long(5420);
	dataBufferOut_long(3483) <= dataBufferIn_long(5421);
	dataBufferOut_long(4226) <= dataBufferIn_long(5422);
	dataBufferOut_long(4969) <= dataBufferIn_long(5423);
	dataBufferOut_long(5712) <= dataBufferIn_long(5424);
	dataBufferOut_long( 311) <= dataBufferIn_long(5425);
	dataBufferOut_long(1054) <= dataBufferIn_long(5426);
	dataBufferOut_long(1797) <= dataBufferIn_long(5427);
	dataBufferOut_long(2540) <= dataBufferIn_long(5428);
	dataBufferOut_long(3283) <= dataBufferIn_long(5429);
	dataBufferOut_long(4026) <= dataBufferIn_long(5430);
	dataBufferOut_long(4769) <= dataBufferIn_long(5431);
	dataBufferOut_long(5512) <= dataBufferIn_long(5432);
	dataBufferOut_long( 111) <= dataBufferIn_long(5433);
	dataBufferOut_long( 854) <= dataBufferIn_long(5434);
	dataBufferOut_long(1597) <= dataBufferIn_long(5435);
	dataBufferOut_long(2340) <= dataBufferIn_long(5436);
	dataBufferOut_long(3083) <= dataBufferIn_long(5437);
	dataBufferOut_long(3826) <= dataBufferIn_long(5438);
	dataBufferOut_long(4569) <= dataBufferIn_long(5439);
	dataBufferOut_long(5312) <= dataBufferIn_long(5440);
	dataBufferOut_long(6055) <= dataBufferIn_long(5441);
	dataBufferOut_long( 654) <= dataBufferIn_long(5442);
	dataBufferOut_long(1397) <= dataBufferIn_long(5443);
	dataBufferOut_long(2140) <= dataBufferIn_long(5444);
	dataBufferOut_long(2883) <= dataBufferIn_long(5445);
	dataBufferOut_long(3626) <= dataBufferIn_long(5446);
	dataBufferOut_long(4369) <= dataBufferIn_long(5447);
	dataBufferOut_long(5112) <= dataBufferIn_long(5448);
	dataBufferOut_long(5855) <= dataBufferIn_long(5449);
	dataBufferOut_long( 454) <= dataBufferIn_long(5450);
	dataBufferOut_long(1197) <= dataBufferIn_long(5451);
	dataBufferOut_long(1940) <= dataBufferIn_long(5452);
	dataBufferOut_long(2683) <= dataBufferIn_long(5453);
	dataBufferOut_long(3426) <= dataBufferIn_long(5454);
	dataBufferOut_long(4169) <= dataBufferIn_long(5455);
	dataBufferOut_long(4912) <= dataBufferIn_long(5456);
	dataBufferOut_long(5655) <= dataBufferIn_long(5457);
	dataBufferOut_long( 254) <= dataBufferIn_long(5458);
	dataBufferOut_long( 997) <= dataBufferIn_long(5459);
	dataBufferOut_long(1740) <= dataBufferIn_long(5460);
	dataBufferOut_long(2483) <= dataBufferIn_long(5461);
	dataBufferOut_long(3226) <= dataBufferIn_long(5462);
	dataBufferOut_long(3969) <= dataBufferIn_long(5463);
	dataBufferOut_long(4712) <= dataBufferIn_long(5464);
	dataBufferOut_long(5455) <= dataBufferIn_long(5465);
	dataBufferOut_long(  54) <= dataBufferIn_long(5466);
	dataBufferOut_long( 797) <= dataBufferIn_long(5467);
	dataBufferOut_long(1540) <= dataBufferIn_long(5468);
	dataBufferOut_long(2283) <= dataBufferIn_long(5469);
	dataBufferOut_long(3026) <= dataBufferIn_long(5470);
	dataBufferOut_long(3769) <= dataBufferIn_long(5471);
	dataBufferOut_long(4512) <= dataBufferIn_long(5472);
	dataBufferOut_long(5255) <= dataBufferIn_long(5473);
	dataBufferOut_long(5998) <= dataBufferIn_long(5474);
	dataBufferOut_long( 597) <= dataBufferIn_long(5475);
	dataBufferOut_long(1340) <= dataBufferIn_long(5476);
	dataBufferOut_long(2083) <= dataBufferIn_long(5477);
	dataBufferOut_long(2826) <= dataBufferIn_long(5478);
	dataBufferOut_long(3569) <= dataBufferIn_long(5479);
	dataBufferOut_long(4312) <= dataBufferIn_long(5480);
	dataBufferOut_long(5055) <= dataBufferIn_long(5481);
	dataBufferOut_long(5798) <= dataBufferIn_long(5482);
	dataBufferOut_long( 397) <= dataBufferIn_long(5483);
	dataBufferOut_long(1140) <= dataBufferIn_long(5484);
	dataBufferOut_long(1883) <= dataBufferIn_long(5485);
	dataBufferOut_long(2626) <= dataBufferIn_long(5486);
	dataBufferOut_long(3369) <= dataBufferIn_long(5487);
	dataBufferOut_long(4112) <= dataBufferIn_long(5488);
	dataBufferOut_long(4855) <= dataBufferIn_long(5489);
	dataBufferOut_long(5598) <= dataBufferIn_long(5490);
	dataBufferOut_long( 197) <= dataBufferIn_long(5491);
	dataBufferOut_long( 940) <= dataBufferIn_long(5492);
	dataBufferOut_long(1683) <= dataBufferIn_long(5493);
	dataBufferOut_long(2426) <= dataBufferIn_long(5494);
	dataBufferOut_long(3169) <= dataBufferIn_long(5495);
	dataBufferOut_long(3912) <= dataBufferIn_long(5496);
	dataBufferOut_long(4655) <= dataBufferIn_long(5497);
	dataBufferOut_long(5398) <= dataBufferIn_long(5498);
	dataBufferOut_long(6141) <= dataBufferIn_long(5499);
	dataBufferOut_long( 740) <= dataBufferIn_long(5500);
	dataBufferOut_long(1483) <= dataBufferIn_long(5501);
	dataBufferOut_long(2226) <= dataBufferIn_long(5502);
	dataBufferOut_long(2969) <= dataBufferIn_long(5503);
	dataBufferOut_long(3712) <= dataBufferIn_long(5504);
	dataBufferOut_long(4455) <= dataBufferIn_long(5505);
	dataBufferOut_long(5198) <= dataBufferIn_long(5506);
	dataBufferOut_long(5941) <= dataBufferIn_long(5507);
	dataBufferOut_long( 540) <= dataBufferIn_long(5508);
	dataBufferOut_long(1283) <= dataBufferIn_long(5509);
	dataBufferOut_long(2026) <= dataBufferIn_long(5510);
	dataBufferOut_long(2769) <= dataBufferIn_long(5511);
	dataBufferOut_long(3512) <= dataBufferIn_long(5512);
	dataBufferOut_long(4255) <= dataBufferIn_long(5513);
	dataBufferOut_long(4998) <= dataBufferIn_long(5514);
	dataBufferOut_long(5741) <= dataBufferIn_long(5515);
	dataBufferOut_long( 340) <= dataBufferIn_long(5516);
	dataBufferOut_long(1083) <= dataBufferIn_long(5517);
	dataBufferOut_long(1826) <= dataBufferIn_long(5518);
	dataBufferOut_long(2569) <= dataBufferIn_long(5519);
	dataBufferOut_long(3312) <= dataBufferIn_long(5520);
	dataBufferOut_long(4055) <= dataBufferIn_long(5521);
	dataBufferOut_long(4798) <= dataBufferIn_long(5522);
	dataBufferOut_long(5541) <= dataBufferIn_long(5523);
	dataBufferOut_long( 140) <= dataBufferIn_long(5524);
	dataBufferOut_long( 883) <= dataBufferIn_long(5525);
	dataBufferOut_long(1626) <= dataBufferIn_long(5526);
	dataBufferOut_long(2369) <= dataBufferIn_long(5527);
	dataBufferOut_long(3112) <= dataBufferIn_long(5528);
	dataBufferOut_long(3855) <= dataBufferIn_long(5529);
	dataBufferOut_long(4598) <= dataBufferIn_long(5530);
	dataBufferOut_long(5341) <= dataBufferIn_long(5531);
	dataBufferOut_long(6084) <= dataBufferIn_long(5532);
	dataBufferOut_long( 683) <= dataBufferIn_long(5533);
	dataBufferOut_long(1426) <= dataBufferIn_long(5534);
	dataBufferOut_long(2169) <= dataBufferIn_long(5535);
	dataBufferOut_long(2912) <= dataBufferIn_long(5536);
	dataBufferOut_long(3655) <= dataBufferIn_long(5537);
	dataBufferOut_long(4398) <= dataBufferIn_long(5538);
	dataBufferOut_long(5141) <= dataBufferIn_long(5539);
	dataBufferOut_long(5884) <= dataBufferIn_long(5540);
	dataBufferOut_long( 483) <= dataBufferIn_long(5541);
	dataBufferOut_long(1226) <= dataBufferIn_long(5542);
	dataBufferOut_long(1969) <= dataBufferIn_long(5543);
	dataBufferOut_long(2712) <= dataBufferIn_long(5544);
	dataBufferOut_long(3455) <= dataBufferIn_long(5545);
	dataBufferOut_long(4198) <= dataBufferIn_long(5546);
	dataBufferOut_long(4941) <= dataBufferIn_long(5547);
	dataBufferOut_long(5684) <= dataBufferIn_long(5548);
	dataBufferOut_long( 283) <= dataBufferIn_long(5549);
	dataBufferOut_long(1026) <= dataBufferIn_long(5550);
	dataBufferOut_long(1769) <= dataBufferIn_long(5551);
	dataBufferOut_long(2512) <= dataBufferIn_long(5552);
	dataBufferOut_long(3255) <= dataBufferIn_long(5553);
	dataBufferOut_long(3998) <= dataBufferIn_long(5554);
	dataBufferOut_long(4741) <= dataBufferIn_long(5555);
	dataBufferOut_long(5484) <= dataBufferIn_long(5556);
	dataBufferOut_long(  83) <= dataBufferIn_long(5557);
	dataBufferOut_long( 826) <= dataBufferIn_long(5558);
	dataBufferOut_long(1569) <= dataBufferIn_long(5559);
	dataBufferOut_long(2312) <= dataBufferIn_long(5560);
	dataBufferOut_long(3055) <= dataBufferIn_long(5561);
	dataBufferOut_long(3798) <= dataBufferIn_long(5562);
	dataBufferOut_long(4541) <= dataBufferIn_long(5563);
	dataBufferOut_long(5284) <= dataBufferIn_long(5564);
	dataBufferOut_long(6027) <= dataBufferIn_long(5565);
	dataBufferOut_long( 626) <= dataBufferIn_long(5566);
	dataBufferOut_long(1369) <= dataBufferIn_long(5567);
	dataBufferOut_long(2112) <= dataBufferIn_long(5568);
	dataBufferOut_long(2855) <= dataBufferIn_long(5569);
	dataBufferOut_long(3598) <= dataBufferIn_long(5570);
	dataBufferOut_long(4341) <= dataBufferIn_long(5571);
	dataBufferOut_long(5084) <= dataBufferIn_long(5572);
	dataBufferOut_long(5827) <= dataBufferIn_long(5573);
	dataBufferOut_long( 426) <= dataBufferIn_long(5574);
	dataBufferOut_long(1169) <= dataBufferIn_long(5575);
	dataBufferOut_long(1912) <= dataBufferIn_long(5576);
	dataBufferOut_long(2655) <= dataBufferIn_long(5577);
	dataBufferOut_long(3398) <= dataBufferIn_long(5578);
	dataBufferOut_long(4141) <= dataBufferIn_long(5579);
	dataBufferOut_long(4884) <= dataBufferIn_long(5580);
	dataBufferOut_long(5627) <= dataBufferIn_long(5581);
	dataBufferOut_long( 226) <= dataBufferIn_long(5582);
	dataBufferOut_long( 969) <= dataBufferIn_long(5583);
	dataBufferOut_long(1712) <= dataBufferIn_long(5584);
	dataBufferOut_long(2455) <= dataBufferIn_long(5585);
	dataBufferOut_long(3198) <= dataBufferIn_long(5586);
	dataBufferOut_long(3941) <= dataBufferIn_long(5587);
	dataBufferOut_long(4684) <= dataBufferIn_long(5588);
	dataBufferOut_long(5427) <= dataBufferIn_long(5589);
	dataBufferOut_long(  26) <= dataBufferIn_long(5590);
	dataBufferOut_long( 769) <= dataBufferIn_long(5591);
	dataBufferOut_long(1512) <= dataBufferIn_long(5592);
	dataBufferOut_long(2255) <= dataBufferIn_long(5593);
	dataBufferOut_long(2998) <= dataBufferIn_long(5594);
	dataBufferOut_long(3741) <= dataBufferIn_long(5595);
	dataBufferOut_long(4484) <= dataBufferIn_long(5596);
	dataBufferOut_long(5227) <= dataBufferIn_long(5597);
	dataBufferOut_long(5970) <= dataBufferIn_long(5598);
	dataBufferOut_long( 569) <= dataBufferIn_long(5599);
	dataBufferOut_long(1312) <= dataBufferIn_long(5600);
	dataBufferOut_long(2055) <= dataBufferIn_long(5601);
	dataBufferOut_long(2798) <= dataBufferIn_long(5602);
	dataBufferOut_long(3541) <= dataBufferIn_long(5603);
	dataBufferOut_long(4284) <= dataBufferIn_long(5604);
	dataBufferOut_long(5027) <= dataBufferIn_long(5605);
	dataBufferOut_long(5770) <= dataBufferIn_long(5606);
	dataBufferOut_long( 369) <= dataBufferIn_long(5607);
	dataBufferOut_long(1112) <= dataBufferIn_long(5608);
	dataBufferOut_long(1855) <= dataBufferIn_long(5609);
	dataBufferOut_long(2598) <= dataBufferIn_long(5610);
	dataBufferOut_long(3341) <= dataBufferIn_long(5611);
	dataBufferOut_long(4084) <= dataBufferIn_long(5612);
	dataBufferOut_long(4827) <= dataBufferIn_long(5613);
	dataBufferOut_long(5570) <= dataBufferIn_long(5614);
	dataBufferOut_long( 169) <= dataBufferIn_long(5615);
	dataBufferOut_long( 912) <= dataBufferIn_long(5616);
	dataBufferOut_long(1655) <= dataBufferIn_long(5617);
	dataBufferOut_long(2398) <= dataBufferIn_long(5618);
	dataBufferOut_long(3141) <= dataBufferIn_long(5619);
	dataBufferOut_long(3884) <= dataBufferIn_long(5620);
	dataBufferOut_long(4627) <= dataBufferIn_long(5621);
	dataBufferOut_long(5370) <= dataBufferIn_long(5622);
	dataBufferOut_long(6113) <= dataBufferIn_long(5623);
	dataBufferOut_long( 712) <= dataBufferIn_long(5624);
	dataBufferOut_long(1455) <= dataBufferIn_long(5625);
	dataBufferOut_long(2198) <= dataBufferIn_long(5626);
	dataBufferOut_long(2941) <= dataBufferIn_long(5627);
	dataBufferOut_long(3684) <= dataBufferIn_long(5628);
	dataBufferOut_long(4427) <= dataBufferIn_long(5629);
	dataBufferOut_long(5170) <= dataBufferIn_long(5630);
	dataBufferOut_long(5913) <= dataBufferIn_long(5631);
	dataBufferOut_long( 512) <= dataBufferIn_long(5632);
	dataBufferOut_long(1255) <= dataBufferIn_long(5633);
	dataBufferOut_long(1998) <= dataBufferIn_long(5634);
	dataBufferOut_long(2741) <= dataBufferIn_long(5635);
	dataBufferOut_long(3484) <= dataBufferIn_long(5636);
	dataBufferOut_long(4227) <= dataBufferIn_long(5637);
	dataBufferOut_long(4970) <= dataBufferIn_long(5638);
	dataBufferOut_long(5713) <= dataBufferIn_long(5639);
	dataBufferOut_long( 312) <= dataBufferIn_long(5640);
	dataBufferOut_long(1055) <= dataBufferIn_long(5641);
	dataBufferOut_long(1798) <= dataBufferIn_long(5642);
	dataBufferOut_long(2541) <= dataBufferIn_long(5643);
	dataBufferOut_long(3284) <= dataBufferIn_long(5644);
	dataBufferOut_long(4027) <= dataBufferIn_long(5645);
	dataBufferOut_long(4770) <= dataBufferIn_long(5646);
	dataBufferOut_long(5513) <= dataBufferIn_long(5647);
	dataBufferOut_long( 112) <= dataBufferIn_long(5648);
	dataBufferOut_long( 855) <= dataBufferIn_long(5649);
	dataBufferOut_long(1598) <= dataBufferIn_long(5650);
	dataBufferOut_long(2341) <= dataBufferIn_long(5651);
	dataBufferOut_long(3084) <= dataBufferIn_long(5652);
	dataBufferOut_long(3827) <= dataBufferIn_long(5653);
	dataBufferOut_long(4570) <= dataBufferIn_long(5654);
	dataBufferOut_long(5313) <= dataBufferIn_long(5655);
	dataBufferOut_long(6056) <= dataBufferIn_long(5656);
	dataBufferOut_long( 655) <= dataBufferIn_long(5657);
	dataBufferOut_long(1398) <= dataBufferIn_long(5658);
	dataBufferOut_long(2141) <= dataBufferIn_long(5659);
	dataBufferOut_long(2884) <= dataBufferIn_long(5660);
	dataBufferOut_long(3627) <= dataBufferIn_long(5661);
	dataBufferOut_long(4370) <= dataBufferIn_long(5662);
	dataBufferOut_long(5113) <= dataBufferIn_long(5663);
	dataBufferOut_long(5856) <= dataBufferIn_long(5664);
	dataBufferOut_long( 455) <= dataBufferIn_long(5665);
	dataBufferOut_long(1198) <= dataBufferIn_long(5666);
	dataBufferOut_long(1941) <= dataBufferIn_long(5667);
	dataBufferOut_long(2684) <= dataBufferIn_long(5668);
	dataBufferOut_long(3427) <= dataBufferIn_long(5669);
	dataBufferOut_long(4170) <= dataBufferIn_long(5670);
	dataBufferOut_long(4913) <= dataBufferIn_long(5671);
	dataBufferOut_long(5656) <= dataBufferIn_long(5672);
	dataBufferOut_long( 255) <= dataBufferIn_long(5673);
	dataBufferOut_long( 998) <= dataBufferIn_long(5674);
	dataBufferOut_long(1741) <= dataBufferIn_long(5675);
	dataBufferOut_long(2484) <= dataBufferIn_long(5676);
	dataBufferOut_long(3227) <= dataBufferIn_long(5677);
	dataBufferOut_long(3970) <= dataBufferIn_long(5678);
	dataBufferOut_long(4713) <= dataBufferIn_long(5679);
	dataBufferOut_long(5456) <= dataBufferIn_long(5680);
	dataBufferOut_long(  55) <= dataBufferIn_long(5681);
	dataBufferOut_long( 798) <= dataBufferIn_long(5682);
	dataBufferOut_long(1541) <= dataBufferIn_long(5683);
	dataBufferOut_long(2284) <= dataBufferIn_long(5684);
	dataBufferOut_long(3027) <= dataBufferIn_long(5685);
	dataBufferOut_long(3770) <= dataBufferIn_long(5686);
	dataBufferOut_long(4513) <= dataBufferIn_long(5687);
	dataBufferOut_long(5256) <= dataBufferIn_long(5688);
	dataBufferOut_long(5999) <= dataBufferIn_long(5689);
	dataBufferOut_long( 598) <= dataBufferIn_long(5690);
	dataBufferOut_long(1341) <= dataBufferIn_long(5691);
	dataBufferOut_long(2084) <= dataBufferIn_long(5692);
	dataBufferOut_long(2827) <= dataBufferIn_long(5693);
	dataBufferOut_long(3570) <= dataBufferIn_long(5694);
	dataBufferOut_long(4313) <= dataBufferIn_long(5695);
	dataBufferOut_long(5056) <= dataBufferIn_long(5696);
	dataBufferOut_long(5799) <= dataBufferIn_long(5697);
	dataBufferOut_long( 398) <= dataBufferIn_long(5698);
	dataBufferOut_long(1141) <= dataBufferIn_long(5699);
	dataBufferOut_long(1884) <= dataBufferIn_long(5700);
	dataBufferOut_long(2627) <= dataBufferIn_long(5701);
	dataBufferOut_long(3370) <= dataBufferIn_long(5702);
	dataBufferOut_long(4113) <= dataBufferIn_long(5703);
	dataBufferOut_long(4856) <= dataBufferIn_long(5704);
	dataBufferOut_long(5599) <= dataBufferIn_long(5705);
	dataBufferOut_long( 198) <= dataBufferIn_long(5706);
	dataBufferOut_long( 941) <= dataBufferIn_long(5707);
	dataBufferOut_long(1684) <= dataBufferIn_long(5708);
	dataBufferOut_long(2427) <= dataBufferIn_long(5709);
	dataBufferOut_long(3170) <= dataBufferIn_long(5710);
	dataBufferOut_long(3913) <= dataBufferIn_long(5711);
	dataBufferOut_long(4656) <= dataBufferIn_long(5712);
	dataBufferOut_long(5399) <= dataBufferIn_long(5713);
	dataBufferOut_long(6142) <= dataBufferIn_long(5714);
	dataBufferOut_long( 741) <= dataBufferIn_long(5715);
	dataBufferOut_long(1484) <= dataBufferIn_long(5716);
	dataBufferOut_long(2227) <= dataBufferIn_long(5717);
	dataBufferOut_long(2970) <= dataBufferIn_long(5718);
	dataBufferOut_long(3713) <= dataBufferIn_long(5719);
	dataBufferOut_long(4456) <= dataBufferIn_long(5720);
	dataBufferOut_long(5199) <= dataBufferIn_long(5721);
	dataBufferOut_long(5942) <= dataBufferIn_long(5722);
	dataBufferOut_long( 541) <= dataBufferIn_long(5723);
	dataBufferOut_long(1284) <= dataBufferIn_long(5724);
	dataBufferOut_long(2027) <= dataBufferIn_long(5725);
	dataBufferOut_long(2770) <= dataBufferIn_long(5726);
	dataBufferOut_long(3513) <= dataBufferIn_long(5727);
	dataBufferOut_long(4256) <= dataBufferIn_long(5728);
	dataBufferOut_long(4999) <= dataBufferIn_long(5729);
	dataBufferOut_long(5742) <= dataBufferIn_long(5730);
	dataBufferOut_long( 341) <= dataBufferIn_long(5731);
	dataBufferOut_long(1084) <= dataBufferIn_long(5732);
	dataBufferOut_long(1827) <= dataBufferIn_long(5733);
	dataBufferOut_long(2570) <= dataBufferIn_long(5734);
	dataBufferOut_long(3313) <= dataBufferIn_long(5735);
	dataBufferOut_long(4056) <= dataBufferIn_long(5736);
	dataBufferOut_long(4799) <= dataBufferIn_long(5737);
	dataBufferOut_long(5542) <= dataBufferIn_long(5738);
	dataBufferOut_long( 141) <= dataBufferIn_long(5739);
	dataBufferOut_long( 884) <= dataBufferIn_long(5740);
	dataBufferOut_long(1627) <= dataBufferIn_long(5741);
	dataBufferOut_long(2370) <= dataBufferIn_long(5742);
	dataBufferOut_long(3113) <= dataBufferIn_long(5743);
	dataBufferOut_long(3856) <= dataBufferIn_long(5744);
	dataBufferOut_long(4599) <= dataBufferIn_long(5745);
	dataBufferOut_long(5342) <= dataBufferIn_long(5746);
	dataBufferOut_long(6085) <= dataBufferIn_long(5747);
	dataBufferOut_long( 684) <= dataBufferIn_long(5748);
	dataBufferOut_long(1427) <= dataBufferIn_long(5749);
	dataBufferOut_long(2170) <= dataBufferIn_long(5750);
	dataBufferOut_long(2913) <= dataBufferIn_long(5751);
	dataBufferOut_long(3656) <= dataBufferIn_long(5752);
	dataBufferOut_long(4399) <= dataBufferIn_long(5753);
	dataBufferOut_long(5142) <= dataBufferIn_long(5754);
	dataBufferOut_long(5885) <= dataBufferIn_long(5755);
	dataBufferOut_long( 484) <= dataBufferIn_long(5756);
	dataBufferOut_long(1227) <= dataBufferIn_long(5757);
	dataBufferOut_long(1970) <= dataBufferIn_long(5758);
	dataBufferOut_long(2713) <= dataBufferIn_long(5759);
	dataBufferOut_long(3456) <= dataBufferIn_long(5760);
	dataBufferOut_long(4199) <= dataBufferIn_long(5761);
	dataBufferOut_long(4942) <= dataBufferIn_long(5762);
	dataBufferOut_long(5685) <= dataBufferIn_long(5763);
	dataBufferOut_long( 284) <= dataBufferIn_long(5764);
	dataBufferOut_long(1027) <= dataBufferIn_long(5765);
	dataBufferOut_long(1770) <= dataBufferIn_long(5766);
	dataBufferOut_long(2513) <= dataBufferIn_long(5767);
	dataBufferOut_long(3256) <= dataBufferIn_long(5768);
	dataBufferOut_long(3999) <= dataBufferIn_long(5769);
	dataBufferOut_long(4742) <= dataBufferIn_long(5770);
	dataBufferOut_long(5485) <= dataBufferIn_long(5771);
	dataBufferOut_long(  84) <= dataBufferIn_long(5772);
	dataBufferOut_long( 827) <= dataBufferIn_long(5773);
	dataBufferOut_long(1570) <= dataBufferIn_long(5774);
	dataBufferOut_long(2313) <= dataBufferIn_long(5775);
	dataBufferOut_long(3056) <= dataBufferIn_long(5776);
	dataBufferOut_long(3799) <= dataBufferIn_long(5777);
	dataBufferOut_long(4542) <= dataBufferIn_long(5778);
	dataBufferOut_long(5285) <= dataBufferIn_long(5779);
	dataBufferOut_long(6028) <= dataBufferIn_long(5780);
	dataBufferOut_long( 627) <= dataBufferIn_long(5781);
	dataBufferOut_long(1370) <= dataBufferIn_long(5782);
	dataBufferOut_long(2113) <= dataBufferIn_long(5783);
	dataBufferOut_long(2856) <= dataBufferIn_long(5784);
	dataBufferOut_long(3599) <= dataBufferIn_long(5785);
	dataBufferOut_long(4342) <= dataBufferIn_long(5786);
	dataBufferOut_long(5085) <= dataBufferIn_long(5787);
	dataBufferOut_long(5828) <= dataBufferIn_long(5788);
	dataBufferOut_long( 427) <= dataBufferIn_long(5789);
	dataBufferOut_long(1170) <= dataBufferIn_long(5790);
	dataBufferOut_long(1913) <= dataBufferIn_long(5791);
	dataBufferOut_long(2656) <= dataBufferIn_long(5792);
	dataBufferOut_long(3399) <= dataBufferIn_long(5793);
	dataBufferOut_long(4142) <= dataBufferIn_long(5794);
	dataBufferOut_long(4885) <= dataBufferIn_long(5795);
	dataBufferOut_long(5628) <= dataBufferIn_long(5796);
	dataBufferOut_long( 227) <= dataBufferIn_long(5797);
	dataBufferOut_long( 970) <= dataBufferIn_long(5798);
	dataBufferOut_long(1713) <= dataBufferIn_long(5799);
	dataBufferOut_long(2456) <= dataBufferIn_long(5800);
	dataBufferOut_long(3199) <= dataBufferIn_long(5801);
	dataBufferOut_long(3942) <= dataBufferIn_long(5802);
	dataBufferOut_long(4685) <= dataBufferIn_long(5803);
	dataBufferOut_long(5428) <= dataBufferIn_long(5804);
	dataBufferOut_long(  27) <= dataBufferIn_long(5805);
	dataBufferOut_long( 770) <= dataBufferIn_long(5806);
	dataBufferOut_long(1513) <= dataBufferIn_long(5807);
	dataBufferOut_long(2256) <= dataBufferIn_long(5808);
	dataBufferOut_long(2999) <= dataBufferIn_long(5809);
	dataBufferOut_long(3742) <= dataBufferIn_long(5810);
	dataBufferOut_long(4485) <= dataBufferIn_long(5811);
	dataBufferOut_long(5228) <= dataBufferIn_long(5812);
	dataBufferOut_long(5971) <= dataBufferIn_long(5813);
	dataBufferOut_long( 570) <= dataBufferIn_long(5814);
	dataBufferOut_long(1313) <= dataBufferIn_long(5815);
	dataBufferOut_long(2056) <= dataBufferIn_long(5816);
	dataBufferOut_long(2799) <= dataBufferIn_long(5817);
	dataBufferOut_long(3542) <= dataBufferIn_long(5818);
	dataBufferOut_long(4285) <= dataBufferIn_long(5819);
	dataBufferOut_long(5028) <= dataBufferIn_long(5820);
	dataBufferOut_long(5771) <= dataBufferIn_long(5821);
	dataBufferOut_long( 370) <= dataBufferIn_long(5822);
	dataBufferOut_long(1113) <= dataBufferIn_long(5823);
	dataBufferOut_long(1856) <= dataBufferIn_long(5824);
	dataBufferOut_long(2599) <= dataBufferIn_long(5825);
	dataBufferOut_long(3342) <= dataBufferIn_long(5826);
	dataBufferOut_long(4085) <= dataBufferIn_long(5827);
	dataBufferOut_long(4828) <= dataBufferIn_long(5828);
	dataBufferOut_long(5571) <= dataBufferIn_long(5829);
	dataBufferOut_long( 170) <= dataBufferIn_long(5830);
	dataBufferOut_long( 913) <= dataBufferIn_long(5831);
	dataBufferOut_long(1656) <= dataBufferIn_long(5832);
	dataBufferOut_long(2399) <= dataBufferIn_long(5833);
	dataBufferOut_long(3142) <= dataBufferIn_long(5834);
	dataBufferOut_long(3885) <= dataBufferIn_long(5835);
	dataBufferOut_long(4628) <= dataBufferIn_long(5836);
	dataBufferOut_long(5371) <= dataBufferIn_long(5837);
	dataBufferOut_long(6114) <= dataBufferIn_long(5838);
	dataBufferOut_long( 713) <= dataBufferIn_long(5839);
	dataBufferOut_long(1456) <= dataBufferIn_long(5840);
	dataBufferOut_long(2199) <= dataBufferIn_long(5841);
	dataBufferOut_long(2942) <= dataBufferIn_long(5842);
	dataBufferOut_long(3685) <= dataBufferIn_long(5843);
	dataBufferOut_long(4428) <= dataBufferIn_long(5844);
	dataBufferOut_long(5171) <= dataBufferIn_long(5845);
	dataBufferOut_long(5914) <= dataBufferIn_long(5846);
	dataBufferOut_long( 513) <= dataBufferIn_long(5847);
	dataBufferOut_long(1256) <= dataBufferIn_long(5848);
	dataBufferOut_long(1999) <= dataBufferIn_long(5849);
	dataBufferOut_long(2742) <= dataBufferIn_long(5850);
	dataBufferOut_long(3485) <= dataBufferIn_long(5851);
	dataBufferOut_long(4228) <= dataBufferIn_long(5852);
	dataBufferOut_long(4971) <= dataBufferIn_long(5853);
	dataBufferOut_long(5714) <= dataBufferIn_long(5854);
	dataBufferOut_long( 313) <= dataBufferIn_long(5855);
	dataBufferOut_long(1056) <= dataBufferIn_long(5856);
	dataBufferOut_long(1799) <= dataBufferIn_long(5857);
	dataBufferOut_long(2542) <= dataBufferIn_long(5858);
	dataBufferOut_long(3285) <= dataBufferIn_long(5859);
	dataBufferOut_long(4028) <= dataBufferIn_long(5860);
	dataBufferOut_long(4771) <= dataBufferIn_long(5861);
	dataBufferOut_long(5514) <= dataBufferIn_long(5862);
	dataBufferOut_long( 113) <= dataBufferIn_long(5863);
	dataBufferOut_long( 856) <= dataBufferIn_long(5864);
	dataBufferOut_long(1599) <= dataBufferIn_long(5865);
	dataBufferOut_long(2342) <= dataBufferIn_long(5866);
	dataBufferOut_long(3085) <= dataBufferIn_long(5867);
	dataBufferOut_long(3828) <= dataBufferIn_long(5868);
	dataBufferOut_long(4571) <= dataBufferIn_long(5869);
	dataBufferOut_long(5314) <= dataBufferIn_long(5870);
	dataBufferOut_long(6057) <= dataBufferIn_long(5871);
	dataBufferOut_long( 656) <= dataBufferIn_long(5872);
	dataBufferOut_long(1399) <= dataBufferIn_long(5873);
	dataBufferOut_long(2142) <= dataBufferIn_long(5874);
	dataBufferOut_long(2885) <= dataBufferIn_long(5875);
	dataBufferOut_long(3628) <= dataBufferIn_long(5876);
	dataBufferOut_long(4371) <= dataBufferIn_long(5877);
	dataBufferOut_long(5114) <= dataBufferIn_long(5878);
	dataBufferOut_long(5857) <= dataBufferIn_long(5879);
	dataBufferOut_long( 456) <= dataBufferIn_long(5880);
	dataBufferOut_long(1199) <= dataBufferIn_long(5881);
	dataBufferOut_long(1942) <= dataBufferIn_long(5882);
	dataBufferOut_long(2685) <= dataBufferIn_long(5883);
	dataBufferOut_long(3428) <= dataBufferIn_long(5884);
	dataBufferOut_long(4171) <= dataBufferIn_long(5885);
	dataBufferOut_long(4914) <= dataBufferIn_long(5886);
	dataBufferOut_long(5657) <= dataBufferIn_long(5887);
	dataBufferOut_long( 256) <= dataBufferIn_long(5888);
	dataBufferOut_long( 999) <= dataBufferIn_long(5889);
	dataBufferOut_long(1742) <= dataBufferIn_long(5890);
	dataBufferOut_long(2485) <= dataBufferIn_long(5891);
	dataBufferOut_long(3228) <= dataBufferIn_long(5892);
	dataBufferOut_long(3971) <= dataBufferIn_long(5893);
	dataBufferOut_long(4714) <= dataBufferIn_long(5894);
	dataBufferOut_long(5457) <= dataBufferIn_long(5895);
	dataBufferOut_long(  56) <= dataBufferIn_long(5896);
	dataBufferOut_long( 799) <= dataBufferIn_long(5897);
	dataBufferOut_long(1542) <= dataBufferIn_long(5898);
	dataBufferOut_long(2285) <= dataBufferIn_long(5899);
	dataBufferOut_long(3028) <= dataBufferIn_long(5900);
	dataBufferOut_long(3771) <= dataBufferIn_long(5901);
	dataBufferOut_long(4514) <= dataBufferIn_long(5902);
	dataBufferOut_long(5257) <= dataBufferIn_long(5903);
	dataBufferOut_long(6000) <= dataBufferIn_long(5904);
	dataBufferOut_long( 599) <= dataBufferIn_long(5905);
	dataBufferOut_long(1342) <= dataBufferIn_long(5906);
	dataBufferOut_long(2085) <= dataBufferIn_long(5907);
	dataBufferOut_long(2828) <= dataBufferIn_long(5908);
	dataBufferOut_long(3571) <= dataBufferIn_long(5909);
	dataBufferOut_long(4314) <= dataBufferIn_long(5910);
	dataBufferOut_long(5057) <= dataBufferIn_long(5911);
	dataBufferOut_long(5800) <= dataBufferIn_long(5912);
	dataBufferOut_long( 399) <= dataBufferIn_long(5913);
	dataBufferOut_long(1142) <= dataBufferIn_long(5914);
	dataBufferOut_long(1885) <= dataBufferIn_long(5915);
	dataBufferOut_long(2628) <= dataBufferIn_long(5916);
	dataBufferOut_long(3371) <= dataBufferIn_long(5917);
	dataBufferOut_long(4114) <= dataBufferIn_long(5918);
	dataBufferOut_long(4857) <= dataBufferIn_long(5919);
	dataBufferOut_long(5600) <= dataBufferIn_long(5920);
	dataBufferOut_long( 199) <= dataBufferIn_long(5921);
	dataBufferOut_long( 942) <= dataBufferIn_long(5922);
	dataBufferOut_long(1685) <= dataBufferIn_long(5923);
	dataBufferOut_long(2428) <= dataBufferIn_long(5924);
	dataBufferOut_long(3171) <= dataBufferIn_long(5925);
	dataBufferOut_long(3914) <= dataBufferIn_long(5926);
	dataBufferOut_long(4657) <= dataBufferIn_long(5927);
	dataBufferOut_long(5400) <= dataBufferIn_long(5928);
	dataBufferOut_long(6143) <= dataBufferIn_long(5929);
	dataBufferOut_long( 742) <= dataBufferIn_long(5930);
	dataBufferOut_long(1485) <= dataBufferIn_long(5931);
	dataBufferOut_long(2228) <= dataBufferIn_long(5932);
	dataBufferOut_long(2971) <= dataBufferIn_long(5933);
	dataBufferOut_long(3714) <= dataBufferIn_long(5934);
	dataBufferOut_long(4457) <= dataBufferIn_long(5935);
	dataBufferOut_long(5200) <= dataBufferIn_long(5936);
	dataBufferOut_long(5943) <= dataBufferIn_long(5937);
	dataBufferOut_long( 542) <= dataBufferIn_long(5938);
	dataBufferOut_long(1285) <= dataBufferIn_long(5939);
	dataBufferOut_long(2028) <= dataBufferIn_long(5940);
	dataBufferOut_long(2771) <= dataBufferIn_long(5941);
	dataBufferOut_long(3514) <= dataBufferIn_long(5942);
	dataBufferOut_long(4257) <= dataBufferIn_long(5943);
	dataBufferOut_long(5000) <= dataBufferIn_long(5944);
	dataBufferOut_long(5743) <= dataBufferIn_long(5945);
	dataBufferOut_long( 342) <= dataBufferIn_long(5946);
	dataBufferOut_long(1085) <= dataBufferIn_long(5947);
	dataBufferOut_long(1828) <= dataBufferIn_long(5948);
	dataBufferOut_long(2571) <= dataBufferIn_long(5949);
	dataBufferOut_long(3314) <= dataBufferIn_long(5950);
	dataBufferOut_long(4057) <= dataBufferIn_long(5951);
	dataBufferOut_long(4800) <= dataBufferIn_long(5952);
	dataBufferOut_long(5543) <= dataBufferIn_long(5953);
	dataBufferOut_long( 142) <= dataBufferIn_long(5954);
	dataBufferOut_long( 885) <= dataBufferIn_long(5955);
	dataBufferOut_long(1628) <= dataBufferIn_long(5956);
	dataBufferOut_long(2371) <= dataBufferIn_long(5957);
	dataBufferOut_long(3114) <= dataBufferIn_long(5958);
	dataBufferOut_long(3857) <= dataBufferIn_long(5959);
	dataBufferOut_long(4600) <= dataBufferIn_long(5960);
	dataBufferOut_long(5343) <= dataBufferIn_long(5961);
	dataBufferOut_long(6086) <= dataBufferIn_long(5962);
	dataBufferOut_long( 685) <= dataBufferIn_long(5963);
	dataBufferOut_long(1428) <= dataBufferIn_long(5964);
	dataBufferOut_long(2171) <= dataBufferIn_long(5965);
	dataBufferOut_long(2914) <= dataBufferIn_long(5966);
	dataBufferOut_long(3657) <= dataBufferIn_long(5967);
	dataBufferOut_long(4400) <= dataBufferIn_long(5968);
	dataBufferOut_long(5143) <= dataBufferIn_long(5969);
	dataBufferOut_long(5886) <= dataBufferIn_long(5970);
	dataBufferOut_long( 485) <= dataBufferIn_long(5971);
	dataBufferOut_long(1228) <= dataBufferIn_long(5972);
	dataBufferOut_long(1971) <= dataBufferIn_long(5973);
	dataBufferOut_long(2714) <= dataBufferIn_long(5974);
	dataBufferOut_long(3457) <= dataBufferIn_long(5975);
	dataBufferOut_long(4200) <= dataBufferIn_long(5976);
	dataBufferOut_long(4943) <= dataBufferIn_long(5977);
	dataBufferOut_long(5686) <= dataBufferIn_long(5978);
	dataBufferOut_long( 285) <= dataBufferIn_long(5979);
	dataBufferOut_long(1028) <= dataBufferIn_long(5980);
	dataBufferOut_long(1771) <= dataBufferIn_long(5981);
	dataBufferOut_long(2514) <= dataBufferIn_long(5982);
	dataBufferOut_long(3257) <= dataBufferIn_long(5983);
	dataBufferOut_long(4000) <= dataBufferIn_long(5984);
	dataBufferOut_long(4743) <= dataBufferIn_long(5985);
	dataBufferOut_long(5486) <= dataBufferIn_long(5986);
	dataBufferOut_long(  85) <= dataBufferIn_long(5987);
	dataBufferOut_long( 828) <= dataBufferIn_long(5988);
	dataBufferOut_long(1571) <= dataBufferIn_long(5989);
	dataBufferOut_long(2314) <= dataBufferIn_long(5990);
	dataBufferOut_long(3057) <= dataBufferIn_long(5991);
	dataBufferOut_long(3800) <= dataBufferIn_long(5992);
	dataBufferOut_long(4543) <= dataBufferIn_long(5993);
	dataBufferOut_long(5286) <= dataBufferIn_long(5994);
	dataBufferOut_long(6029) <= dataBufferIn_long(5995);
	dataBufferOut_long( 628) <= dataBufferIn_long(5996);
	dataBufferOut_long(1371) <= dataBufferIn_long(5997);
	dataBufferOut_long(2114) <= dataBufferIn_long(5998);
	dataBufferOut_long(2857) <= dataBufferIn_long(5999);
	dataBufferOut_long(3600) <= dataBufferIn_long(6000);
	dataBufferOut_long(4343) <= dataBufferIn_long(6001);
	dataBufferOut_long(5086) <= dataBufferIn_long(6002);
	dataBufferOut_long(5829) <= dataBufferIn_long(6003);
	dataBufferOut_long( 428) <= dataBufferIn_long(6004);
	dataBufferOut_long(1171) <= dataBufferIn_long(6005);
	dataBufferOut_long(1914) <= dataBufferIn_long(6006);
	dataBufferOut_long(2657) <= dataBufferIn_long(6007);
	dataBufferOut_long(3400) <= dataBufferIn_long(6008);
	dataBufferOut_long(4143) <= dataBufferIn_long(6009);
	dataBufferOut_long(4886) <= dataBufferIn_long(6010);
	dataBufferOut_long(5629) <= dataBufferIn_long(6011);
	dataBufferOut_long( 228) <= dataBufferIn_long(6012);
	dataBufferOut_long( 971) <= dataBufferIn_long(6013);
	dataBufferOut_long(1714) <= dataBufferIn_long(6014);
	dataBufferOut_long(2457) <= dataBufferIn_long(6015);
	dataBufferOut_long(3200) <= dataBufferIn_long(6016);
	dataBufferOut_long(3943) <= dataBufferIn_long(6017);
	dataBufferOut_long(4686) <= dataBufferIn_long(6018);
	dataBufferOut_long(5429) <= dataBufferIn_long(6019);
	dataBufferOut_long(  28) <= dataBufferIn_long(6020);
	dataBufferOut_long( 771) <= dataBufferIn_long(6021);
	dataBufferOut_long(1514) <= dataBufferIn_long(6022);
	dataBufferOut_long(2257) <= dataBufferIn_long(6023);
	dataBufferOut_long(3000) <= dataBufferIn_long(6024);
	dataBufferOut_long(3743) <= dataBufferIn_long(6025);
	dataBufferOut_long(4486) <= dataBufferIn_long(6026);
	dataBufferOut_long(5229) <= dataBufferIn_long(6027);
	dataBufferOut_long(5972) <= dataBufferIn_long(6028);
	dataBufferOut_long( 571) <= dataBufferIn_long(6029);
	dataBufferOut_long(1314) <= dataBufferIn_long(6030);
	dataBufferOut_long(2057) <= dataBufferIn_long(6031);
	dataBufferOut_long(2800) <= dataBufferIn_long(6032);
	dataBufferOut_long(3543) <= dataBufferIn_long(6033);
	dataBufferOut_long(4286) <= dataBufferIn_long(6034);
	dataBufferOut_long(5029) <= dataBufferIn_long(6035);
	dataBufferOut_long(5772) <= dataBufferIn_long(6036);
	dataBufferOut_long( 371) <= dataBufferIn_long(6037);
	dataBufferOut_long(1114) <= dataBufferIn_long(6038);
	dataBufferOut_long(1857) <= dataBufferIn_long(6039);
	dataBufferOut_long(2600) <= dataBufferIn_long(6040);
	dataBufferOut_long(3343) <= dataBufferIn_long(6041);
	dataBufferOut_long(4086) <= dataBufferIn_long(6042);
	dataBufferOut_long(4829) <= dataBufferIn_long(6043);
	dataBufferOut_long(5572) <= dataBufferIn_long(6044);
	dataBufferOut_long( 171) <= dataBufferIn_long(6045);
	dataBufferOut_long( 914) <= dataBufferIn_long(6046);
	dataBufferOut_long(1657) <= dataBufferIn_long(6047);
	dataBufferOut_long(2400) <= dataBufferIn_long(6048);
	dataBufferOut_long(3143) <= dataBufferIn_long(6049);
	dataBufferOut_long(3886) <= dataBufferIn_long(6050);
	dataBufferOut_long(4629) <= dataBufferIn_long(6051);
	dataBufferOut_long(5372) <= dataBufferIn_long(6052);
	dataBufferOut_long(6115) <= dataBufferIn_long(6053);
	dataBufferOut_long( 714) <= dataBufferIn_long(6054);
	dataBufferOut_long(1457) <= dataBufferIn_long(6055);
	dataBufferOut_long(2200) <= dataBufferIn_long(6056);
	dataBufferOut_long(2943) <= dataBufferIn_long(6057);
	dataBufferOut_long(3686) <= dataBufferIn_long(6058);
	dataBufferOut_long(4429) <= dataBufferIn_long(6059);
	dataBufferOut_long(5172) <= dataBufferIn_long(6060);
	dataBufferOut_long(5915) <= dataBufferIn_long(6061);
	dataBufferOut_long( 514) <= dataBufferIn_long(6062);
	dataBufferOut_long(1257) <= dataBufferIn_long(6063);
	dataBufferOut_long(2000) <= dataBufferIn_long(6064);
	dataBufferOut_long(2743) <= dataBufferIn_long(6065);
	dataBufferOut_long(3486) <= dataBufferIn_long(6066);
	dataBufferOut_long(4229) <= dataBufferIn_long(6067);
	dataBufferOut_long(4972) <= dataBufferIn_long(6068);
	dataBufferOut_long(5715) <= dataBufferIn_long(6069);
	dataBufferOut_long( 314) <= dataBufferIn_long(6070);
	dataBufferOut_long(1057) <= dataBufferIn_long(6071);
	dataBufferOut_long(1800) <= dataBufferIn_long(6072);
	dataBufferOut_long(2543) <= dataBufferIn_long(6073);
	dataBufferOut_long(3286) <= dataBufferIn_long(6074);
	dataBufferOut_long(4029) <= dataBufferIn_long(6075);
	dataBufferOut_long(4772) <= dataBufferIn_long(6076);
	dataBufferOut_long(5515) <= dataBufferIn_long(6077);
	dataBufferOut_long( 114) <= dataBufferIn_long(6078);
	dataBufferOut_long( 857) <= dataBufferIn_long(6079);
	dataBufferOut_long(1600) <= dataBufferIn_long(6080);
	dataBufferOut_long(2343) <= dataBufferIn_long(6081);
	dataBufferOut_long(3086) <= dataBufferIn_long(6082);
	dataBufferOut_long(3829) <= dataBufferIn_long(6083);
	dataBufferOut_long(4572) <= dataBufferIn_long(6084);
	dataBufferOut_long(5315) <= dataBufferIn_long(6085);
	dataBufferOut_long(6058) <= dataBufferIn_long(6086);
	dataBufferOut_long( 657) <= dataBufferIn_long(6087);
	dataBufferOut_long(1400) <= dataBufferIn_long(6088);
	dataBufferOut_long(2143) <= dataBufferIn_long(6089);
	dataBufferOut_long(2886) <= dataBufferIn_long(6090);
	dataBufferOut_long(3629) <= dataBufferIn_long(6091);
	dataBufferOut_long(4372) <= dataBufferIn_long(6092);
	dataBufferOut_long(5115) <= dataBufferIn_long(6093);
	dataBufferOut_long(5858) <= dataBufferIn_long(6094);
	dataBufferOut_long( 457) <= dataBufferIn_long(6095);
	dataBufferOut_long(1200) <= dataBufferIn_long(6096);
	dataBufferOut_long(1943) <= dataBufferIn_long(6097);
	dataBufferOut_long(2686) <= dataBufferIn_long(6098);
	dataBufferOut_long(3429) <= dataBufferIn_long(6099);
	dataBufferOut_long(4172) <= dataBufferIn_long(6100);
	dataBufferOut_long(4915) <= dataBufferIn_long(6101);
	dataBufferOut_long(5658) <= dataBufferIn_long(6102);
	dataBufferOut_long( 257) <= dataBufferIn_long(6103);
	dataBufferOut_long(1000) <= dataBufferIn_long(6104);
	dataBufferOut_long(1743) <= dataBufferIn_long(6105);
	dataBufferOut_long(2486) <= dataBufferIn_long(6106);
	dataBufferOut_long(3229) <= dataBufferIn_long(6107);
	dataBufferOut_long(3972) <= dataBufferIn_long(6108);
	dataBufferOut_long(4715) <= dataBufferIn_long(6109);
	dataBufferOut_long(5458) <= dataBufferIn_long(6110);
	dataBufferOut_long(  57) <= dataBufferIn_long(6111);
	dataBufferOut_long( 800) <= dataBufferIn_long(6112);
	dataBufferOut_long(1543) <= dataBufferIn_long(6113);
	dataBufferOut_long(2286) <= dataBufferIn_long(6114);
	dataBufferOut_long(3029) <= dataBufferIn_long(6115);
	dataBufferOut_long(3772) <= dataBufferIn_long(6116);
	dataBufferOut_long(4515) <= dataBufferIn_long(6117);
	dataBufferOut_long(5258) <= dataBufferIn_long(6118);
	dataBufferOut_long(6001) <= dataBufferIn_long(6119);
	dataBufferOut_long( 600) <= dataBufferIn_long(6120);
	dataBufferOut_long(1343) <= dataBufferIn_long(6121);
	dataBufferOut_long(2086) <= dataBufferIn_long(6122);
	dataBufferOut_long(2829) <= dataBufferIn_long(6123);
	dataBufferOut_long(3572) <= dataBufferIn_long(6124);
	dataBufferOut_long(4315) <= dataBufferIn_long(6125);
	dataBufferOut_long(5058) <= dataBufferIn_long(6126);
	dataBufferOut_long(5801) <= dataBufferIn_long(6127);
	dataBufferOut_long( 400) <= dataBufferIn_long(6128);
	dataBufferOut_long(1143) <= dataBufferIn_long(6129);
	dataBufferOut_long(1886) <= dataBufferIn_long(6130);
	dataBufferOut_long(2629) <= dataBufferIn_long(6131);
	dataBufferOut_long(3372) <= dataBufferIn_long(6132);
	dataBufferOut_long(4115) <= dataBufferIn_long(6133);
	dataBufferOut_long(4858) <= dataBufferIn_long(6134);
	dataBufferOut_long(5601) <= dataBufferIn_long(6135);
	dataBufferOut_long( 200) <= dataBufferIn_long(6136);
	dataBufferOut_long( 943) <= dataBufferIn_long(6137);
	dataBufferOut_long(1686) <= dataBufferIn_long(6138);
	dataBufferOut_long(2429) <= dataBufferIn_long(6139);
	dataBufferOut_long(3172) <= dataBufferIn_long(6140);
	dataBufferOut_long(3915) <= dataBufferIn_long(6141);
	dataBufferOut_long(4658) <= dataBufferIn_long(6142);
	dataBufferOut_long(5401) <= dataBufferIn_long(6143);


end arch1;


library ieee;
use ieee.std_logic_1164.all;

entity TurboInterleaver_Interleaver is
	port (
		clk, reset_async:			in std_logic;
		flag_long:					in std_logic;

		dataBufferIn:			in std_logic_vector(6143 DOWNTO 0);
		dataBufferOut:			out std_logic_vector(6143 DOWNTO 0)
	);
end TurboInterleaver_Interleaver;

architecture arch1 of TurboInterleaver_Interleaver is

begin

	dataBufferOut(   0) <= dataBufferIn(   0) when (flag_long='1') else '0';
	dataBufferOut(   1) <= dataBufferIn( 743) when (flag_long='1') else '0';
	dataBufferOut(   2) <= dataBufferIn(1486) when (flag_long='1') else '0';
	dataBufferOut(   3) <= dataBufferIn(2229) when (flag_long='1') else '0';
	dataBufferOut(   4) <= dataBufferIn(2972) when (flag_long='1') else '0';
	dataBufferOut(   5) <= dataBufferIn(3715) when (flag_long='1') else '0';
	dataBufferOut(   6) <= dataBufferIn(4458) when (flag_long='1') else '0';
	dataBufferOut(   7) <= dataBufferIn(5201) when (flag_long='1') else '0';
	dataBufferOut(   8) <= dataBufferIn(5944) when (flag_long='1') else '0';
	dataBufferOut(   9) <= dataBufferIn( 543) when (flag_long='1') else '0';
	dataBufferOut(  10) <= dataBufferIn(1286) when (flag_long='1') else '0';
	dataBufferOut(  11) <= dataBufferIn(2029) when (flag_long='1') else '0';
	dataBufferOut(  12) <= dataBufferIn(2772) when (flag_long='1') else '0';
	dataBufferOut(  13) <= dataBufferIn(3515) when (flag_long='1') else '0';
	dataBufferOut(  14) <= dataBufferIn(4258) when (flag_long='1') else '0';
	dataBufferOut(  15) <= dataBufferIn(5001) when (flag_long='1') else '0';
	dataBufferOut(  16) <= dataBufferIn(5744) when (flag_long='1') else '0';
	dataBufferOut(  17) <= dataBufferIn( 343) when (flag_long='1') else '0';
	dataBufferOut(  18) <= dataBufferIn(1086) when (flag_long='1') else '0';
	dataBufferOut(  19) <= dataBufferIn(1829) when (flag_long='1') else '0';
	dataBufferOut(  20) <= dataBufferIn(2572) when (flag_long='1') else '0';
	dataBufferOut(  21) <= dataBufferIn(3315) when (flag_long='1') else '0';
	dataBufferOut(  22) <= dataBufferIn(4058) when (flag_long='1') else '0';
	dataBufferOut(  23) <= dataBufferIn(4801) when (flag_long='1') else '0';
	dataBufferOut(  24) <= dataBufferIn(5544) when (flag_long='1') else '0';
	dataBufferOut(  25) <= dataBufferIn( 143) when (flag_long='1') else '0';
	dataBufferOut(  26) <= dataBufferIn( 886) when (flag_long='1') else '0';
	dataBufferOut(  27) <= dataBufferIn(1629) when (flag_long='1') else '0';
	dataBufferOut(  28) <= dataBufferIn(2372) when (flag_long='1') else '0';
	dataBufferOut(  29) <= dataBufferIn(3115) when (flag_long='1') else '0';
	dataBufferOut(  30) <= dataBufferIn(3858) when (flag_long='1') else '0';
	dataBufferOut(  31) <= dataBufferIn(4601) when (flag_long='1') else '0';
	dataBufferOut(  32) <= dataBufferIn(5344) when (flag_long='1') else '0';
	dataBufferOut(  33) <= dataBufferIn(6087) when (flag_long='1') else '0';
	dataBufferOut(  34) <= dataBufferIn( 686) when (flag_long='1') else '0';
	dataBufferOut(  35) <= dataBufferIn(1429) when (flag_long='1') else '0';
	dataBufferOut(  36) <= dataBufferIn(2172) when (flag_long='1') else '0';
	dataBufferOut(  37) <= dataBufferIn(2915) when (flag_long='1') else '0';
	dataBufferOut(  38) <= dataBufferIn(3658) when (flag_long='1') else '0';
	dataBufferOut(  39) <= dataBufferIn(4401) when (flag_long='1') else '0';
	dataBufferOut(  40) <= dataBufferIn(5144) when (flag_long='1') else '0';
	dataBufferOut(  41) <= dataBufferIn(5887) when (flag_long='1') else '0';
	dataBufferOut(  42) <= dataBufferIn( 486) when (flag_long='1') else '0';
	dataBufferOut(  43) <= dataBufferIn(1229) when (flag_long='1') else '0';
	dataBufferOut(  44) <= dataBufferIn(1972) when (flag_long='1') else '0';
	dataBufferOut(  45) <= dataBufferIn(2715) when (flag_long='1') else '0';
	dataBufferOut(  46) <= dataBufferIn(3458) when (flag_long='1') else '0';
	dataBufferOut(  47) <= dataBufferIn(4201) when (flag_long='1') else '0';
	dataBufferOut(  48) <= dataBufferIn(4944) when (flag_long='1') else '0';
	dataBufferOut(  49) <= dataBufferIn(5687) when (flag_long='1') else '0';
	dataBufferOut(  50) <= dataBufferIn( 286) when (flag_long='1') else '0';
	dataBufferOut(  51) <= dataBufferIn(1029) when (flag_long='1') else '0';
	dataBufferOut(  52) <= dataBufferIn(1772) when (flag_long='1') else '0';
	dataBufferOut(  53) <= dataBufferIn(2515) when (flag_long='1') else '0';
	dataBufferOut(  54) <= dataBufferIn(3258) when (flag_long='1') else '0';
	dataBufferOut(  55) <= dataBufferIn(4001) when (flag_long='1') else '0';
	dataBufferOut(  56) <= dataBufferIn(4744) when (flag_long='1') else '0';
	dataBufferOut(  57) <= dataBufferIn(5487) when (flag_long='1') else '0';
	dataBufferOut(  58) <= dataBufferIn(  86) when (flag_long='1') else '0';
	dataBufferOut(  59) <= dataBufferIn( 829) when (flag_long='1') else '0';
	dataBufferOut(  60) <= dataBufferIn(1572) when (flag_long='1') else '0';
	dataBufferOut(  61) <= dataBufferIn(2315) when (flag_long='1') else '0';
	dataBufferOut(  62) <= dataBufferIn(3058) when (flag_long='1') else '0';
	dataBufferOut(  63) <= dataBufferIn(3801) when (flag_long='1') else '0';
	dataBufferOut(  64) <= dataBufferIn(4544) when (flag_long='1') else '0';
	dataBufferOut(  65) <= dataBufferIn(5287) when (flag_long='1') else '0';
	dataBufferOut(  66) <= dataBufferIn(6030) when (flag_long='1') else '0';
	dataBufferOut(  67) <= dataBufferIn( 629) when (flag_long='1') else '0';
	dataBufferOut(  68) <= dataBufferIn(1372) when (flag_long='1') else '0';
	dataBufferOut(  69) <= dataBufferIn(2115) when (flag_long='1') else '0';
	dataBufferOut(  70) <= dataBufferIn(2858) when (flag_long='1') else '0';
	dataBufferOut(  71) <= dataBufferIn(3601) when (flag_long='1') else '0';
	dataBufferOut(  72) <= dataBufferIn(4344) when (flag_long='1') else '0';
	dataBufferOut(  73) <= dataBufferIn(5087) when (flag_long='1') else '0';
	dataBufferOut(  74) <= dataBufferIn(5830) when (flag_long='1') else '0';
	dataBufferOut(  75) <= dataBufferIn( 429) when (flag_long='1') else '0';
	dataBufferOut(  76) <= dataBufferIn(1172) when (flag_long='1') else '0';
	dataBufferOut(  77) <= dataBufferIn(1915) when (flag_long='1') else '0';
	dataBufferOut(  78) <= dataBufferIn(2658) when (flag_long='1') else '0';
	dataBufferOut(  79) <= dataBufferIn(3401) when (flag_long='1') else '0';
	dataBufferOut(  80) <= dataBufferIn(4144) when (flag_long='1') else '0';
	dataBufferOut(  81) <= dataBufferIn(4887) when (flag_long='1') else '0';
	dataBufferOut(  82) <= dataBufferIn(5630) when (flag_long='1') else '0';
	dataBufferOut(  83) <= dataBufferIn( 229) when (flag_long='1') else '0';
	dataBufferOut(  84) <= dataBufferIn( 972) when (flag_long='1') else '0';
	dataBufferOut(  85) <= dataBufferIn(1715) when (flag_long='1') else '0';
	dataBufferOut(  86) <= dataBufferIn(2458) when (flag_long='1') else '0';
	dataBufferOut(  87) <= dataBufferIn(3201) when (flag_long='1') else '0';
	dataBufferOut(  88) <= dataBufferIn(3944) when (flag_long='1') else '0';
	dataBufferOut(  89) <= dataBufferIn(4687) when (flag_long='1') else '0';
	dataBufferOut(  90) <= dataBufferIn(5430) when (flag_long='1') else '0';
	dataBufferOut(  91) <= dataBufferIn(  29) when (flag_long='1') else '0';
	dataBufferOut(  92) <= dataBufferIn( 772) when (flag_long='1') else '0';
	dataBufferOut(  93) <= dataBufferIn(1515) when (flag_long='1') else '0';
	dataBufferOut(  94) <= dataBufferIn(2258) when (flag_long='1') else '0';
	dataBufferOut(  95) <= dataBufferIn(3001) when (flag_long='1') else '0';
	dataBufferOut(  96) <= dataBufferIn(3744) when (flag_long='1') else '0';
	dataBufferOut(  97) <= dataBufferIn(4487) when (flag_long='1') else '0';
	dataBufferOut(  98) <= dataBufferIn(5230) when (flag_long='1') else '0';
	dataBufferOut(  99) <= dataBufferIn(5973) when (flag_long='1') else '0';
	dataBufferOut( 100) <= dataBufferIn( 572) when (flag_long='1') else '0';
	dataBufferOut( 101) <= dataBufferIn(1315) when (flag_long='1') else '0';
	dataBufferOut( 102) <= dataBufferIn(2058) when (flag_long='1') else '0';
	dataBufferOut( 103) <= dataBufferIn(2801) when (flag_long='1') else '0';
	dataBufferOut( 104) <= dataBufferIn(3544) when (flag_long='1') else '0';
	dataBufferOut( 105) <= dataBufferIn(4287) when (flag_long='1') else '0';
	dataBufferOut( 106) <= dataBufferIn(5030) when (flag_long='1') else '0';
	dataBufferOut( 107) <= dataBufferIn(5773) when (flag_long='1') else '0';
	dataBufferOut( 108) <= dataBufferIn( 372) when (flag_long='1') else '0';
	dataBufferOut( 109) <= dataBufferIn(1115) when (flag_long='1') else '0';
	dataBufferOut( 110) <= dataBufferIn(1858) when (flag_long='1') else '0';
	dataBufferOut( 111) <= dataBufferIn(2601) when (flag_long='1') else '0';
	dataBufferOut( 112) <= dataBufferIn(3344) when (flag_long='1') else '0';
	dataBufferOut( 113) <= dataBufferIn(4087) when (flag_long='1') else '0';
	dataBufferOut( 114) <= dataBufferIn(4830) when (flag_long='1') else '0';
	dataBufferOut( 115) <= dataBufferIn(5573) when (flag_long='1') else '0';
	dataBufferOut( 116) <= dataBufferIn( 172) when (flag_long='1') else '0';
	dataBufferOut( 117) <= dataBufferIn( 915) when (flag_long='1') else '0';
	dataBufferOut( 118) <= dataBufferIn(1658) when (flag_long='1') else '0';
	dataBufferOut( 119) <= dataBufferIn(2401) when (flag_long='1') else '0';
	dataBufferOut( 120) <= dataBufferIn(3144) when (flag_long='1') else '0';
	dataBufferOut( 121) <= dataBufferIn(3887) when (flag_long='1') else '0';
	dataBufferOut( 122) <= dataBufferIn(4630) when (flag_long='1') else '0';
	dataBufferOut( 123) <= dataBufferIn(5373) when (flag_long='1') else '0';
	dataBufferOut( 124) <= dataBufferIn(6116) when (flag_long='1') else '0';
	dataBufferOut( 125) <= dataBufferIn( 715) when (flag_long='1') else '0';
	dataBufferOut( 126) <= dataBufferIn(1458) when (flag_long='1') else '0';
	dataBufferOut( 127) <= dataBufferIn(2201) when (flag_long='1') else '0';
	dataBufferOut( 128) <= dataBufferIn(2944) when (flag_long='1') else '0';
	dataBufferOut( 129) <= dataBufferIn(3687) when (flag_long='1') else '0';
	dataBufferOut( 130) <= dataBufferIn(4430) when (flag_long='1') else '0';
	dataBufferOut( 131) <= dataBufferIn(5173) when (flag_long='1') else '0';
	dataBufferOut( 132) <= dataBufferIn(5916) when (flag_long='1') else '0';
	dataBufferOut( 133) <= dataBufferIn( 515) when (flag_long='1') else '0';
	dataBufferOut( 134) <= dataBufferIn(1258) when (flag_long='1') else '0';
	dataBufferOut( 135) <= dataBufferIn(2001) when (flag_long='1') else '0';
	dataBufferOut( 136) <= dataBufferIn(2744) when (flag_long='1') else '0';
	dataBufferOut( 137) <= dataBufferIn(3487) when (flag_long='1') else '0';
	dataBufferOut( 138) <= dataBufferIn(4230) when (flag_long='1') else '0';
	dataBufferOut( 139) <= dataBufferIn(4973) when (flag_long='1') else '0';
	dataBufferOut( 140) <= dataBufferIn(5716) when (flag_long='1') else '0';
	dataBufferOut( 141) <= dataBufferIn( 315) when (flag_long='1') else '0';
	dataBufferOut( 142) <= dataBufferIn(1058) when (flag_long='1') else '0';
	dataBufferOut( 143) <= dataBufferIn(1801) when (flag_long='1') else '0';
	dataBufferOut( 144) <= dataBufferIn(2544) when (flag_long='1') else '0';
	dataBufferOut( 145) <= dataBufferIn(3287) when (flag_long='1') else '0';
	dataBufferOut( 146) <= dataBufferIn(4030) when (flag_long='1') else '0';
	dataBufferOut( 147) <= dataBufferIn(4773) when (flag_long='1') else '0';
	dataBufferOut( 148) <= dataBufferIn(5516) when (flag_long='1') else '0';
	dataBufferOut( 149) <= dataBufferIn( 115) when (flag_long='1') else '0';
	dataBufferOut( 150) <= dataBufferIn( 858) when (flag_long='1') else '0';
	dataBufferOut( 151) <= dataBufferIn(1601) when (flag_long='1') else '0';
	dataBufferOut( 152) <= dataBufferIn(2344) when (flag_long='1') else '0';
	dataBufferOut( 153) <= dataBufferIn(3087) when (flag_long='1') else '0';
	dataBufferOut( 154) <= dataBufferIn(3830) when (flag_long='1') else '0';
	dataBufferOut( 155) <= dataBufferIn(4573) when (flag_long='1') else '0';
	dataBufferOut( 156) <= dataBufferIn(5316) when (flag_long='1') else '0';
	dataBufferOut( 157) <= dataBufferIn(6059) when (flag_long='1') else '0';
	dataBufferOut( 158) <= dataBufferIn( 658) when (flag_long='1') else '0';
	dataBufferOut( 159) <= dataBufferIn(1401) when (flag_long='1') else '0';
	dataBufferOut( 160) <= dataBufferIn(2144) when (flag_long='1') else '0';
	dataBufferOut( 161) <= dataBufferIn(2887) when (flag_long='1') else '0';
	dataBufferOut( 162) <= dataBufferIn(3630) when (flag_long='1') else '0';
	dataBufferOut( 163) <= dataBufferIn(4373) when (flag_long='1') else '0';
	dataBufferOut( 164) <= dataBufferIn(5116) when (flag_long='1') else '0';
	dataBufferOut( 165) <= dataBufferIn(5859) when (flag_long='1') else '0';
	dataBufferOut( 166) <= dataBufferIn( 458) when (flag_long='1') else '0';
	dataBufferOut( 167) <= dataBufferIn(1201) when (flag_long='1') else '0';
	dataBufferOut( 168) <= dataBufferIn(1944) when (flag_long='1') else '0';
	dataBufferOut( 169) <= dataBufferIn(2687) when (flag_long='1') else '0';
	dataBufferOut( 170) <= dataBufferIn(3430) when (flag_long='1') else '0';
	dataBufferOut( 171) <= dataBufferIn(4173) when (flag_long='1') else '0';
	dataBufferOut( 172) <= dataBufferIn(4916) when (flag_long='1') else '0';
	dataBufferOut( 173) <= dataBufferIn(5659) when (flag_long='1') else '0';
	dataBufferOut( 174) <= dataBufferIn( 258) when (flag_long='1') else '0';
	dataBufferOut( 175) <= dataBufferIn(1001) when (flag_long='1') else '0';
	dataBufferOut( 176) <= dataBufferIn(1744) when (flag_long='1') else '0';
	dataBufferOut( 177) <= dataBufferIn(2487) when (flag_long='1') else '0';
	dataBufferOut( 178) <= dataBufferIn(3230) when (flag_long='1') else '0';
	dataBufferOut( 179) <= dataBufferIn(3973) when (flag_long='1') else '0';
	dataBufferOut( 180) <= dataBufferIn(4716) when (flag_long='1') else '0';
	dataBufferOut( 181) <= dataBufferIn(5459) when (flag_long='1') else '0';
	dataBufferOut( 182) <= dataBufferIn(  58) when (flag_long='1') else '0';
	dataBufferOut( 183) <= dataBufferIn( 801) when (flag_long='1') else '0';
	dataBufferOut( 184) <= dataBufferIn(1544) when (flag_long='1') else '0';
	dataBufferOut( 185) <= dataBufferIn(2287) when (flag_long='1') else '0';
	dataBufferOut( 186) <= dataBufferIn(3030) when (flag_long='1') else '0';
	dataBufferOut( 187) <= dataBufferIn(3773) when (flag_long='1') else '0';
	dataBufferOut( 188) <= dataBufferIn(4516) when (flag_long='1') else '0';
	dataBufferOut( 189) <= dataBufferIn(5259) when (flag_long='1') else '0';
	dataBufferOut( 190) <= dataBufferIn(6002) when (flag_long='1') else '0';
	dataBufferOut( 191) <= dataBufferIn( 601) when (flag_long='1') else '0';
	dataBufferOut( 192) <= dataBufferIn(1344) when (flag_long='1') else '0';
	dataBufferOut( 193) <= dataBufferIn(2087) when (flag_long='1') else '0';
	dataBufferOut( 194) <= dataBufferIn(2830) when (flag_long='1') else '0';
	dataBufferOut( 195) <= dataBufferIn(3573) when (flag_long='1') else '0';
	dataBufferOut( 196) <= dataBufferIn(4316) when (flag_long='1') else '0';
	dataBufferOut( 197) <= dataBufferIn(5059) when (flag_long='1') else '0';
	dataBufferOut( 198) <= dataBufferIn(5802) when (flag_long='1') else '0';
	dataBufferOut( 199) <= dataBufferIn( 401) when (flag_long='1') else '0';
	dataBufferOut( 200) <= dataBufferIn(1144) when (flag_long='1') else '0';
	dataBufferOut( 201) <= dataBufferIn(1887) when (flag_long='1') else '0';
	dataBufferOut( 202) <= dataBufferIn(2630) when (flag_long='1') else '0';
	dataBufferOut( 203) <= dataBufferIn(3373) when (flag_long='1') else '0';
	dataBufferOut( 204) <= dataBufferIn(4116) when (flag_long='1') else '0';
	dataBufferOut( 205) <= dataBufferIn(4859) when (flag_long='1') else '0';
	dataBufferOut( 206) <= dataBufferIn(5602) when (flag_long='1') else '0';
	dataBufferOut( 207) <= dataBufferIn( 201) when (flag_long='1') else '0';
	dataBufferOut( 208) <= dataBufferIn( 944) when (flag_long='1') else '0';
	dataBufferOut( 209) <= dataBufferIn(1687) when (flag_long='1') else '0';
	dataBufferOut( 210) <= dataBufferIn(2430) when (flag_long='1') else '0';
	dataBufferOut( 211) <= dataBufferIn(3173) when (flag_long='1') else '0';
	dataBufferOut( 212) <= dataBufferIn(3916) when (flag_long='1') else '0';
	dataBufferOut( 213) <= dataBufferIn(4659) when (flag_long='1') else '0';
	dataBufferOut( 214) <= dataBufferIn(5402) when (flag_long='1') else '0';
	dataBufferOut( 215) <= dataBufferIn(   1) when (flag_long='1') else '0';
	dataBufferOut( 216) <= dataBufferIn( 744) when (flag_long='1') else '0';
	dataBufferOut( 217) <= dataBufferIn(1487) when (flag_long='1') else '0';
	dataBufferOut( 218) <= dataBufferIn(2230) when (flag_long='1') else '0';
	dataBufferOut( 219) <= dataBufferIn(2973) when (flag_long='1') else '0';
	dataBufferOut( 220) <= dataBufferIn(3716) when (flag_long='1') else '0';
	dataBufferOut( 221) <= dataBufferIn(4459) when (flag_long='1') else '0';
	dataBufferOut( 222) <= dataBufferIn(5202) when (flag_long='1') else '0';
	dataBufferOut( 223) <= dataBufferIn(5945) when (flag_long='1') else '0';
	dataBufferOut( 224) <= dataBufferIn( 544) when (flag_long='1') else '0';
	dataBufferOut( 225) <= dataBufferIn(1287) when (flag_long='1') else '0';
	dataBufferOut( 226) <= dataBufferIn(2030) when (flag_long='1') else '0';
	dataBufferOut( 227) <= dataBufferIn(2773) when (flag_long='1') else '0';
	dataBufferOut( 228) <= dataBufferIn(3516) when (flag_long='1') else '0';
	dataBufferOut( 229) <= dataBufferIn(4259) when (flag_long='1') else '0';
	dataBufferOut( 230) <= dataBufferIn(5002) when (flag_long='1') else '0';
	dataBufferOut( 231) <= dataBufferIn(5745) when (flag_long='1') else '0';
	dataBufferOut( 232) <= dataBufferIn( 344) when (flag_long='1') else '0';
	dataBufferOut( 233) <= dataBufferIn(1087) when (flag_long='1') else '0';
	dataBufferOut( 234) <= dataBufferIn(1830) when (flag_long='1') else '0';
	dataBufferOut( 235) <= dataBufferIn(2573) when (flag_long='1') else '0';
	dataBufferOut( 236) <= dataBufferIn(3316) when (flag_long='1') else '0';
	dataBufferOut( 237) <= dataBufferIn(4059) when (flag_long='1') else '0';
	dataBufferOut( 238) <= dataBufferIn(4802) when (flag_long='1') else '0';
	dataBufferOut( 239) <= dataBufferIn(5545) when (flag_long='1') else '0';
	dataBufferOut( 240) <= dataBufferIn( 144) when (flag_long='1') else '0';
	dataBufferOut( 241) <= dataBufferIn( 887) when (flag_long='1') else '0';
	dataBufferOut( 242) <= dataBufferIn(1630) when (flag_long='1') else '0';
	dataBufferOut( 243) <= dataBufferIn(2373) when (flag_long='1') else '0';
	dataBufferOut( 244) <= dataBufferIn(3116) when (flag_long='1') else '0';
	dataBufferOut( 245) <= dataBufferIn(3859) when (flag_long='1') else '0';
	dataBufferOut( 246) <= dataBufferIn(4602) when (flag_long='1') else '0';
	dataBufferOut( 247) <= dataBufferIn(5345) when (flag_long='1') else '0';
	dataBufferOut( 248) <= dataBufferIn(6088) when (flag_long='1') else '0';
	dataBufferOut( 249) <= dataBufferIn( 687) when (flag_long='1') else '0';
	dataBufferOut( 250) <= dataBufferIn(1430) when (flag_long='1') else '0';
	dataBufferOut( 251) <= dataBufferIn(2173) when (flag_long='1') else '0';
	dataBufferOut( 252) <= dataBufferIn(2916) when (flag_long='1') else '0';
	dataBufferOut( 253) <= dataBufferIn(3659) when (flag_long='1') else '0';
	dataBufferOut( 254) <= dataBufferIn(4402) when (flag_long='1') else '0';
	dataBufferOut( 255) <= dataBufferIn(5145) when (flag_long='1') else '0';
	dataBufferOut( 256) <= dataBufferIn(5888) when (flag_long='1') else '0';
	dataBufferOut( 257) <= dataBufferIn( 487) when (flag_long='1') else '0';
	dataBufferOut( 258) <= dataBufferIn(1230) when (flag_long='1') else '0';
	dataBufferOut( 259) <= dataBufferIn(1973) when (flag_long='1') else '0';
	dataBufferOut( 260) <= dataBufferIn(2716) when (flag_long='1') else '0';
	dataBufferOut( 261) <= dataBufferIn(3459) when (flag_long='1') else '0';
	dataBufferOut( 262) <= dataBufferIn(4202) when (flag_long='1') else '0';
	dataBufferOut( 263) <= dataBufferIn(4945) when (flag_long='1') else '0';
	dataBufferOut( 264) <= dataBufferIn(5688) when (flag_long='1') else '0';
	dataBufferOut( 265) <= dataBufferIn( 287) when (flag_long='1') else '0';
	dataBufferOut( 266) <= dataBufferIn(1030) when (flag_long='1') else '0';
	dataBufferOut( 267) <= dataBufferIn(1773) when (flag_long='1') else '0';
	dataBufferOut( 268) <= dataBufferIn(2516) when (flag_long='1') else '0';
	dataBufferOut( 269) <= dataBufferIn(3259) when (flag_long='1') else '0';
	dataBufferOut( 270) <= dataBufferIn(4002) when (flag_long='1') else '0';
	dataBufferOut( 271) <= dataBufferIn(4745) when (flag_long='1') else '0';
	dataBufferOut( 272) <= dataBufferIn(5488) when (flag_long='1') else '0';
	dataBufferOut( 273) <= dataBufferIn(  87) when (flag_long='1') else '0';
	dataBufferOut( 274) <= dataBufferIn( 830) when (flag_long='1') else '0';
	dataBufferOut( 275) <= dataBufferIn(1573) when (flag_long='1') else '0';
	dataBufferOut( 276) <= dataBufferIn(2316) when (flag_long='1') else '0';
	dataBufferOut( 277) <= dataBufferIn(3059) when (flag_long='1') else '0';
	dataBufferOut( 278) <= dataBufferIn(3802) when (flag_long='1') else '0';
	dataBufferOut( 279) <= dataBufferIn(4545) when (flag_long='1') else '0';
	dataBufferOut( 280) <= dataBufferIn(5288) when (flag_long='1') else '0';
	dataBufferOut( 281) <= dataBufferIn(6031) when (flag_long='1') else '0';
	dataBufferOut( 282) <= dataBufferIn( 630) when (flag_long='1') else '0';
	dataBufferOut( 283) <= dataBufferIn(1373) when (flag_long='1') else '0';
	dataBufferOut( 284) <= dataBufferIn(2116) when (flag_long='1') else '0';
	dataBufferOut( 285) <= dataBufferIn(2859) when (flag_long='1') else '0';
	dataBufferOut( 286) <= dataBufferIn(3602) when (flag_long='1') else '0';
	dataBufferOut( 287) <= dataBufferIn(4345) when (flag_long='1') else '0';
	dataBufferOut( 288) <= dataBufferIn(5088) when (flag_long='1') else '0';
	dataBufferOut( 289) <= dataBufferIn(5831) when (flag_long='1') else '0';
	dataBufferOut( 290) <= dataBufferIn( 430) when (flag_long='1') else '0';
	dataBufferOut( 291) <= dataBufferIn(1173) when (flag_long='1') else '0';
	dataBufferOut( 292) <= dataBufferIn(1916) when (flag_long='1') else '0';
	dataBufferOut( 293) <= dataBufferIn(2659) when (flag_long='1') else '0';
	dataBufferOut( 294) <= dataBufferIn(3402) when (flag_long='1') else '0';
	dataBufferOut( 295) <= dataBufferIn(4145) when (flag_long='1') else '0';
	dataBufferOut( 296) <= dataBufferIn(4888) when (flag_long='1') else '0';
	dataBufferOut( 297) <= dataBufferIn(5631) when (flag_long='1') else '0';
	dataBufferOut( 298) <= dataBufferIn( 230) when (flag_long='1') else '0';
	dataBufferOut( 299) <= dataBufferIn( 973) when (flag_long='1') else '0';
	dataBufferOut( 300) <= dataBufferIn(1716) when (flag_long='1') else '0';
	dataBufferOut( 301) <= dataBufferIn(2459) when (flag_long='1') else '0';
	dataBufferOut( 302) <= dataBufferIn(3202) when (flag_long='1') else '0';
	dataBufferOut( 303) <= dataBufferIn(3945) when (flag_long='1') else '0';
	dataBufferOut( 304) <= dataBufferIn(4688) when (flag_long='1') else '0';
	dataBufferOut( 305) <= dataBufferIn(5431) when (flag_long='1') else '0';
	dataBufferOut( 306) <= dataBufferIn(  30) when (flag_long='1') else '0';
	dataBufferOut( 307) <= dataBufferIn( 773) when (flag_long='1') else '0';
	dataBufferOut( 308) <= dataBufferIn(1516) when (flag_long='1') else '0';
	dataBufferOut( 309) <= dataBufferIn(2259) when (flag_long='1') else '0';
	dataBufferOut( 310) <= dataBufferIn(3002) when (flag_long='1') else '0';
	dataBufferOut( 311) <= dataBufferIn(3745) when (flag_long='1') else '0';
	dataBufferOut( 312) <= dataBufferIn(4488) when (flag_long='1') else '0';
	dataBufferOut( 313) <= dataBufferIn(5231) when (flag_long='1') else '0';
	dataBufferOut( 314) <= dataBufferIn(5974) when (flag_long='1') else '0';
	dataBufferOut( 315) <= dataBufferIn( 573) when (flag_long='1') else '0';
	dataBufferOut( 316) <= dataBufferIn(1316) when (flag_long='1') else '0';
	dataBufferOut( 317) <= dataBufferIn(2059) when (flag_long='1') else '0';
	dataBufferOut( 318) <= dataBufferIn(2802) when (flag_long='1') else '0';
	dataBufferOut( 319) <= dataBufferIn(3545) when (flag_long='1') else '0';
	dataBufferOut( 320) <= dataBufferIn(4288) when (flag_long='1') else '0';
	dataBufferOut( 321) <= dataBufferIn(5031) when (flag_long='1') else '0';
	dataBufferOut( 322) <= dataBufferIn(5774) when (flag_long='1') else '0';
	dataBufferOut( 323) <= dataBufferIn( 373) when (flag_long='1') else '0';
	dataBufferOut( 324) <= dataBufferIn(1116) when (flag_long='1') else '0';
	dataBufferOut( 325) <= dataBufferIn(1859) when (flag_long='1') else '0';
	dataBufferOut( 326) <= dataBufferIn(2602) when (flag_long='1') else '0';
	dataBufferOut( 327) <= dataBufferIn(3345) when (flag_long='1') else '0';
	dataBufferOut( 328) <= dataBufferIn(4088) when (flag_long='1') else '0';
	dataBufferOut( 329) <= dataBufferIn(4831) when (flag_long='1') else '0';
	dataBufferOut( 330) <= dataBufferIn(5574) when (flag_long='1') else '0';
	dataBufferOut( 331) <= dataBufferIn( 173) when (flag_long='1') else '0';
	dataBufferOut( 332) <= dataBufferIn( 916) when (flag_long='1') else '0';
	dataBufferOut( 333) <= dataBufferIn(1659) when (flag_long='1') else '0';
	dataBufferOut( 334) <= dataBufferIn(2402) when (flag_long='1') else '0';
	dataBufferOut( 335) <= dataBufferIn(3145) when (flag_long='1') else '0';
	dataBufferOut( 336) <= dataBufferIn(3888) when (flag_long='1') else '0';
	dataBufferOut( 337) <= dataBufferIn(4631) when (flag_long='1') else '0';
	dataBufferOut( 338) <= dataBufferIn(5374) when (flag_long='1') else '0';
	dataBufferOut( 339) <= dataBufferIn(6117) when (flag_long='1') else '0';
	dataBufferOut( 340) <= dataBufferIn( 716) when (flag_long='1') else '0';
	dataBufferOut( 341) <= dataBufferIn(1459) when (flag_long='1') else '0';
	dataBufferOut( 342) <= dataBufferIn(2202) when (flag_long='1') else '0';
	dataBufferOut( 343) <= dataBufferIn(2945) when (flag_long='1') else '0';
	dataBufferOut( 344) <= dataBufferIn(3688) when (flag_long='1') else '0';
	dataBufferOut( 345) <= dataBufferIn(4431) when (flag_long='1') else '0';
	dataBufferOut( 346) <= dataBufferIn(5174) when (flag_long='1') else '0';
	dataBufferOut( 347) <= dataBufferIn(5917) when (flag_long='1') else '0';
	dataBufferOut( 348) <= dataBufferIn( 516) when (flag_long='1') else '0';
	dataBufferOut( 349) <= dataBufferIn(1259) when (flag_long='1') else '0';
	dataBufferOut( 350) <= dataBufferIn(2002) when (flag_long='1') else '0';
	dataBufferOut( 351) <= dataBufferIn(2745) when (flag_long='1') else '0';
	dataBufferOut( 352) <= dataBufferIn(3488) when (flag_long='1') else '0';
	dataBufferOut( 353) <= dataBufferIn(4231) when (flag_long='1') else '0';
	dataBufferOut( 354) <= dataBufferIn(4974) when (flag_long='1') else '0';
	dataBufferOut( 355) <= dataBufferIn(5717) when (flag_long='1') else '0';
	dataBufferOut( 356) <= dataBufferIn( 316) when (flag_long='1') else '0';
	dataBufferOut( 357) <= dataBufferIn(1059) when (flag_long='1') else '0';
	dataBufferOut( 358) <= dataBufferIn(1802) when (flag_long='1') else '0';
	dataBufferOut( 359) <= dataBufferIn(2545) when (flag_long='1') else '0';
	dataBufferOut( 360) <= dataBufferIn(3288) when (flag_long='1') else '0';
	dataBufferOut( 361) <= dataBufferIn(4031) when (flag_long='1') else '0';
	dataBufferOut( 362) <= dataBufferIn(4774) when (flag_long='1') else '0';
	dataBufferOut( 363) <= dataBufferIn(5517) when (flag_long='1') else '0';
	dataBufferOut( 364) <= dataBufferIn( 116) when (flag_long='1') else '0';
	dataBufferOut( 365) <= dataBufferIn( 859) when (flag_long='1') else '0';
	dataBufferOut( 366) <= dataBufferIn(1602) when (flag_long='1') else '0';
	dataBufferOut( 367) <= dataBufferIn(2345) when (flag_long='1') else '0';
	dataBufferOut( 368) <= dataBufferIn(3088) when (flag_long='1') else '0';
	dataBufferOut( 369) <= dataBufferIn(3831) when (flag_long='1') else '0';
	dataBufferOut( 370) <= dataBufferIn(4574) when (flag_long='1') else '0';
	dataBufferOut( 371) <= dataBufferIn(5317) when (flag_long='1') else '0';
	dataBufferOut( 372) <= dataBufferIn(6060) when (flag_long='1') else '0';
	dataBufferOut( 373) <= dataBufferIn( 659) when (flag_long='1') else '0';
	dataBufferOut( 374) <= dataBufferIn(1402) when (flag_long='1') else '0';
	dataBufferOut( 375) <= dataBufferIn(2145) when (flag_long='1') else '0';
	dataBufferOut( 376) <= dataBufferIn(2888) when (flag_long='1') else '0';
	dataBufferOut( 377) <= dataBufferIn(3631) when (flag_long='1') else '0';
	dataBufferOut( 378) <= dataBufferIn(4374) when (flag_long='1') else '0';
	dataBufferOut( 379) <= dataBufferIn(5117) when (flag_long='1') else '0';
	dataBufferOut( 380) <= dataBufferIn(5860) when (flag_long='1') else '0';
	dataBufferOut( 381) <= dataBufferIn( 459) when (flag_long='1') else '0';
	dataBufferOut( 382) <= dataBufferIn(1202) when (flag_long='1') else '0';
	dataBufferOut( 383) <= dataBufferIn(1945) when (flag_long='1') else '0';
	dataBufferOut( 384) <= dataBufferIn(2688) when (flag_long='1') else '0';
	dataBufferOut( 385) <= dataBufferIn(3431) when (flag_long='1') else '0';
	dataBufferOut( 386) <= dataBufferIn(4174) when (flag_long='1') else '0';
	dataBufferOut( 387) <= dataBufferIn(4917) when (flag_long='1') else '0';
	dataBufferOut( 388) <= dataBufferIn(5660) when (flag_long='1') else '0';
	dataBufferOut( 389) <= dataBufferIn( 259) when (flag_long='1') else '0';
	dataBufferOut( 390) <= dataBufferIn(1002) when (flag_long='1') else '0';
	dataBufferOut( 391) <= dataBufferIn(1745) when (flag_long='1') else '0';
	dataBufferOut( 392) <= dataBufferIn(2488) when (flag_long='1') else '0';
	dataBufferOut( 393) <= dataBufferIn(3231) when (flag_long='1') else '0';
	dataBufferOut( 394) <= dataBufferIn(3974) when (flag_long='1') else '0';
	dataBufferOut( 395) <= dataBufferIn(4717) when (flag_long='1') else '0';
	dataBufferOut( 396) <= dataBufferIn(5460) when (flag_long='1') else '0';
	dataBufferOut( 397) <= dataBufferIn(  59) when (flag_long='1') else '0';
	dataBufferOut( 398) <= dataBufferIn( 802) when (flag_long='1') else '0';
	dataBufferOut( 399) <= dataBufferIn(1545) when (flag_long='1') else '0';
	dataBufferOut( 400) <= dataBufferIn(2288) when (flag_long='1') else '0';
	dataBufferOut( 401) <= dataBufferIn(3031) when (flag_long='1') else '0';
	dataBufferOut( 402) <= dataBufferIn(3774) when (flag_long='1') else '0';
	dataBufferOut( 403) <= dataBufferIn(4517) when (flag_long='1') else '0';
	dataBufferOut( 404) <= dataBufferIn(5260) when (flag_long='1') else '0';
	dataBufferOut( 405) <= dataBufferIn(6003) when (flag_long='1') else '0';
	dataBufferOut( 406) <= dataBufferIn( 602) when (flag_long='1') else '0';
	dataBufferOut( 407) <= dataBufferIn(1345) when (flag_long='1') else '0';
	dataBufferOut( 408) <= dataBufferIn(2088) when (flag_long='1') else '0';
	dataBufferOut( 409) <= dataBufferIn(2831) when (flag_long='1') else '0';
	dataBufferOut( 410) <= dataBufferIn(3574) when (flag_long='1') else '0';
	dataBufferOut( 411) <= dataBufferIn(4317) when (flag_long='1') else '0';
	dataBufferOut( 412) <= dataBufferIn(5060) when (flag_long='1') else '0';
	dataBufferOut( 413) <= dataBufferIn(5803) when (flag_long='1') else '0';
	dataBufferOut( 414) <= dataBufferIn( 402) when (flag_long='1') else '0';
	dataBufferOut( 415) <= dataBufferIn(1145) when (flag_long='1') else '0';
	dataBufferOut( 416) <= dataBufferIn(1888) when (flag_long='1') else '0';
	dataBufferOut( 417) <= dataBufferIn(2631) when (flag_long='1') else '0';
	dataBufferOut( 418) <= dataBufferIn(3374) when (flag_long='1') else '0';
	dataBufferOut( 419) <= dataBufferIn(4117) when (flag_long='1') else '0';
	dataBufferOut( 420) <= dataBufferIn(4860) when (flag_long='1') else '0';
	dataBufferOut( 421) <= dataBufferIn(5603) when (flag_long='1') else '0';
	dataBufferOut( 422) <= dataBufferIn( 202) when (flag_long='1') else '0';
	dataBufferOut( 423) <= dataBufferIn( 945) when (flag_long='1') else '0';
	dataBufferOut( 424) <= dataBufferIn(1688) when (flag_long='1') else '0';
	dataBufferOut( 425) <= dataBufferIn(2431) when (flag_long='1') else '0';
	dataBufferOut( 426) <= dataBufferIn(3174) when (flag_long='1') else '0';
	dataBufferOut( 427) <= dataBufferIn(3917) when (flag_long='1') else '0';
	dataBufferOut( 428) <= dataBufferIn(4660) when (flag_long='1') else '0';
	dataBufferOut( 429) <= dataBufferIn(5403) when (flag_long='1') else '0';
	dataBufferOut( 430) <= dataBufferIn(   2) when (flag_long='1') else '0';
	dataBufferOut( 431) <= dataBufferIn( 745) when (flag_long='1') else '0';
	dataBufferOut( 432) <= dataBufferIn(1488) when (flag_long='1') else '0';
	dataBufferOut( 433) <= dataBufferIn(2231) when (flag_long='1') else '0';
	dataBufferOut( 434) <= dataBufferIn(2974) when (flag_long='1') else '0';
	dataBufferOut( 435) <= dataBufferIn(3717) when (flag_long='1') else '0';
	dataBufferOut( 436) <= dataBufferIn(4460) when (flag_long='1') else '0';
	dataBufferOut( 437) <= dataBufferIn(5203) when (flag_long='1') else '0';
	dataBufferOut( 438) <= dataBufferIn(5946) when (flag_long='1') else '0';
	dataBufferOut( 439) <= dataBufferIn( 545) when (flag_long='1') else '0';
	dataBufferOut( 440) <= dataBufferIn(1288) when (flag_long='1') else '0';
	dataBufferOut( 441) <= dataBufferIn(2031) when (flag_long='1') else '0';
	dataBufferOut( 442) <= dataBufferIn(2774) when (flag_long='1') else '0';
	dataBufferOut( 443) <= dataBufferIn(3517) when (flag_long='1') else '0';
	dataBufferOut( 444) <= dataBufferIn(4260) when (flag_long='1') else '0';
	dataBufferOut( 445) <= dataBufferIn(5003) when (flag_long='1') else '0';
	dataBufferOut( 446) <= dataBufferIn(5746) when (flag_long='1') else '0';
	dataBufferOut( 447) <= dataBufferIn( 345) when (flag_long='1') else '0';
	dataBufferOut( 448) <= dataBufferIn(1088) when (flag_long='1') else '0';
	dataBufferOut( 449) <= dataBufferIn(1831) when (flag_long='1') else '0';
	dataBufferOut( 450) <= dataBufferIn(2574) when (flag_long='1') else '0';
	dataBufferOut( 451) <= dataBufferIn(3317) when (flag_long='1') else '0';
	dataBufferOut( 452) <= dataBufferIn(4060) when (flag_long='1') else '0';
	dataBufferOut( 453) <= dataBufferIn(4803) when (flag_long='1') else '0';
	dataBufferOut( 454) <= dataBufferIn(5546) when (flag_long='1') else '0';
	dataBufferOut( 455) <= dataBufferIn( 145) when (flag_long='1') else '0';
	dataBufferOut( 456) <= dataBufferIn( 888) when (flag_long='1') else '0';
	dataBufferOut( 457) <= dataBufferIn(1631) when (flag_long='1') else '0';
	dataBufferOut( 458) <= dataBufferIn(2374) when (flag_long='1') else '0';
	dataBufferOut( 459) <= dataBufferIn(3117) when (flag_long='1') else '0';
	dataBufferOut( 460) <= dataBufferIn(3860) when (flag_long='1') else '0';
	dataBufferOut( 461) <= dataBufferIn(4603) when (flag_long='1') else '0';
	dataBufferOut( 462) <= dataBufferIn(5346) when (flag_long='1') else '0';
	dataBufferOut( 463) <= dataBufferIn(6089) when (flag_long='1') else '0';
	dataBufferOut( 464) <= dataBufferIn( 688) when (flag_long='1') else '0';
	dataBufferOut( 465) <= dataBufferIn(1431) when (flag_long='1') else '0';
	dataBufferOut( 466) <= dataBufferIn(2174) when (flag_long='1') else '0';
	dataBufferOut( 467) <= dataBufferIn(2917) when (flag_long='1') else '0';
	dataBufferOut( 468) <= dataBufferIn(3660) when (flag_long='1') else '0';
	dataBufferOut( 469) <= dataBufferIn(4403) when (flag_long='1') else '0';
	dataBufferOut( 470) <= dataBufferIn(5146) when (flag_long='1') else '0';
	dataBufferOut( 471) <= dataBufferIn(5889) when (flag_long='1') else '0';
	dataBufferOut( 472) <= dataBufferIn( 488) when (flag_long='1') else '0';
	dataBufferOut( 473) <= dataBufferIn(1231) when (flag_long='1') else '0';
	dataBufferOut( 474) <= dataBufferIn(1974) when (flag_long='1') else '0';
	dataBufferOut( 475) <= dataBufferIn(2717) when (flag_long='1') else '0';
	dataBufferOut( 476) <= dataBufferIn(3460) when (flag_long='1') else '0';
	dataBufferOut( 477) <= dataBufferIn(4203) when (flag_long='1') else '0';
	dataBufferOut( 478) <= dataBufferIn(4946) when (flag_long='1') else '0';
	dataBufferOut( 479) <= dataBufferIn(5689) when (flag_long='1') else '0';
	dataBufferOut( 480) <= dataBufferIn( 288) when (flag_long='1') else '0';
	dataBufferOut( 481) <= dataBufferIn(1031) when (flag_long='1') else '0';
	dataBufferOut( 482) <= dataBufferIn(1774) when (flag_long='1') else '0';
	dataBufferOut( 483) <= dataBufferIn(2517) when (flag_long='1') else '0';
	dataBufferOut( 484) <= dataBufferIn(3260) when (flag_long='1') else '0';
	dataBufferOut( 485) <= dataBufferIn(4003) when (flag_long='1') else '0';
	dataBufferOut( 486) <= dataBufferIn(4746) when (flag_long='1') else '0';
	dataBufferOut( 487) <= dataBufferIn(5489) when (flag_long='1') else '0';
	dataBufferOut( 488) <= dataBufferIn(  88) when (flag_long='1') else '0';
	dataBufferOut( 489) <= dataBufferIn( 831) when (flag_long='1') else '0';
	dataBufferOut( 490) <= dataBufferIn(1574) when (flag_long='1') else '0';
	dataBufferOut( 491) <= dataBufferIn(2317) when (flag_long='1') else '0';
	dataBufferOut( 492) <= dataBufferIn(3060) when (flag_long='1') else '0';
	dataBufferOut( 493) <= dataBufferIn(3803) when (flag_long='1') else '0';
	dataBufferOut( 494) <= dataBufferIn(4546) when (flag_long='1') else '0';
	dataBufferOut( 495) <= dataBufferIn(5289) when (flag_long='1') else '0';
	dataBufferOut( 496) <= dataBufferIn(6032) when (flag_long='1') else '0';
	dataBufferOut( 497) <= dataBufferIn( 631) when (flag_long='1') else '0';
	dataBufferOut( 498) <= dataBufferIn(1374) when (flag_long='1') else '0';
	dataBufferOut( 499) <= dataBufferIn(2117) when (flag_long='1') else '0';
	dataBufferOut( 500) <= dataBufferIn(2860) when (flag_long='1') else '0';
	dataBufferOut( 501) <= dataBufferIn(3603) when (flag_long='1') else '0';
	dataBufferOut( 502) <= dataBufferIn(4346) when (flag_long='1') else '0';
	dataBufferOut( 503) <= dataBufferIn(5089) when (flag_long='1') else '0';
	dataBufferOut( 504) <= dataBufferIn(5832) when (flag_long='1') else '0';
	dataBufferOut( 505) <= dataBufferIn( 431) when (flag_long='1') else '0';
	dataBufferOut( 506) <= dataBufferIn(1174) when (flag_long='1') else '0';
	dataBufferOut( 507) <= dataBufferIn(1917) when (flag_long='1') else '0';
	dataBufferOut( 508) <= dataBufferIn(2660) when (flag_long='1') else '0';
	dataBufferOut( 509) <= dataBufferIn(3403) when (flag_long='1') else '0';
	dataBufferOut( 510) <= dataBufferIn(4146) when (flag_long='1') else '0';
	dataBufferOut( 511) <= dataBufferIn(4889) when (flag_long='1') else '0';
	dataBufferOut( 512) <= dataBufferIn(5632) when (flag_long='1') else '0';
	dataBufferOut( 513) <= dataBufferIn( 231) when (flag_long='1') else '0';
	dataBufferOut( 514) <= dataBufferIn( 974) when (flag_long='1') else '0';
	dataBufferOut( 515) <= dataBufferIn(1717) when (flag_long='1') else '0';
	dataBufferOut( 516) <= dataBufferIn(2460) when (flag_long='1') else '0';
	dataBufferOut( 517) <= dataBufferIn(3203) when (flag_long='1') else '0';
	dataBufferOut( 518) <= dataBufferIn(3946) when (flag_long='1') else '0';
	dataBufferOut( 519) <= dataBufferIn(4689) when (flag_long='1') else '0';
	dataBufferOut( 520) <= dataBufferIn(5432) when (flag_long='1') else '0';
	dataBufferOut( 521) <= dataBufferIn(  31) when (flag_long='1') else '0';
	dataBufferOut( 522) <= dataBufferIn( 774) when (flag_long='1') else '0';
	dataBufferOut( 523) <= dataBufferIn(1517) when (flag_long='1') else '0';
	dataBufferOut( 524) <= dataBufferIn(2260) when (flag_long='1') else '0';
	dataBufferOut( 525) <= dataBufferIn(3003) when (flag_long='1') else '0';
	dataBufferOut( 526) <= dataBufferIn(3746) when (flag_long='1') else '0';
	dataBufferOut( 527) <= dataBufferIn(4489) when (flag_long='1') else '0';
	dataBufferOut( 528) <= dataBufferIn(5232) when (flag_long='1') else '0';
	dataBufferOut( 529) <= dataBufferIn(5975) when (flag_long='1') else '0';
	dataBufferOut( 530) <= dataBufferIn( 574) when (flag_long='1') else '0';
	dataBufferOut( 531) <= dataBufferIn(1317) when (flag_long='1') else '0';
	dataBufferOut( 532) <= dataBufferIn(2060) when (flag_long='1') else '0';
	dataBufferOut( 533) <= dataBufferIn(2803) when (flag_long='1') else '0';
	dataBufferOut( 534) <= dataBufferIn(3546) when (flag_long='1') else '0';
	dataBufferOut( 535) <= dataBufferIn(4289) when (flag_long='1') else '0';
	dataBufferOut( 536) <= dataBufferIn(5032) when (flag_long='1') else '0';
	dataBufferOut( 537) <= dataBufferIn(5775) when (flag_long='1') else '0';
	dataBufferOut( 538) <= dataBufferIn( 374) when (flag_long='1') else '0';
	dataBufferOut( 539) <= dataBufferIn(1117) when (flag_long='1') else '0';
	dataBufferOut( 540) <= dataBufferIn(1860) when (flag_long='1') else '0';
	dataBufferOut( 541) <= dataBufferIn(2603) when (flag_long='1') else '0';
	dataBufferOut( 542) <= dataBufferIn(3346) when (flag_long='1') else '0';
	dataBufferOut( 543) <= dataBufferIn(4089) when (flag_long='1') else '0';
	dataBufferOut( 544) <= dataBufferIn(4832) when (flag_long='1') else '0';
	dataBufferOut( 545) <= dataBufferIn(5575) when (flag_long='1') else '0';
	dataBufferOut( 546) <= dataBufferIn( 174) when (flag_long='1') else '0';
	dataBufferOut( 547) <= dataBufferIn( 917) when (flag_long='1') else '0';
	dataBufferOut( 548) <= dataBufferIn(1660) when (flag_long='1') else '0';
	dataBufferOut( 549) <= dataBufferIn(2403) when (flag_long='1') else '0';
	dataBufferOut( 550) <= dataBufferIn(3146) when (flag_long='1') else '0';
	dataBufferOut( 551) <= dataBufferIn(3889) when (flag_long='1') else '0';
	dataBufferOut( 552) <= dataBufferIn(4632) when (flag_long='1') else '0';
	dataBufferOut( 553) <= dataBufferIn(5375) when (flag_long='1') else '0';
	dataBufferOut( 554) <= dataBufferIn(6118) when (flag_long='1') else '0';
	dataBufferOut( 555) <= dataBufferIn( 717) when (flag_long='1') else '0';
	dataBufferOut( 556) <= dataBufferIn(1460) when (flag_long='1') else '0';
	dataBufferOut( 557) <= dataBufferIn(2203) when (flag_long='1') else '0';
	dataBufferOut( 558) <= dataBufferIn(2946) when (flag_long='1') else '0';
	dataBufferOut( 559) <= dataBufferIn(3689) when (flag_long='1') else '0';
	dataBufferOut( 560) <= dataBufferIn(4432) when (flag_long='1') else '0';
	dataBufferOut( 561) <= dataBufferIn(5175) when (flag_long='1') else '0';
	dataBufferOut( 562) <= dataBufferIn(5918) when (flag_long='1') else '0';
	dataBufferOut( 563) <= dataBufferIn( 517) when (flag_long='1') else '0';
	dataBufferOut( 564) <= dataBufferIn(1260) when (flag_long='1') else '0';
	dataBufferOut( 565) <= dataBufferIn(2003) when (flag_long='1') else '0';
	dataBufferOut( 566) <= dataBufferIn(2746) when (flag_long='1') else '0';
	dataBufferOut( 567) <= dataBufferIn(3489) when (flag_long='1') else '0';
	dataBufferOut( 568) <= dataBufferIn(4232) when (flag_long='1') else '0';
	dataBufferOut( 569) <= dataBufferIn(4975) when (flag_long='1') else '0';
	dataBufferOut( 570) <= dataBufferIn(5718) when (flag_long='1') else '0';
	dataBufferOut( 571) <= dataBufferIn( 317) when (flag_long='1') else '0';
	dataBufferOut( 572) <= dataBufferIn(1060) when (flag_long='1') else '0';
	dataBufferOut( 573) <= dataBufferIn(1803) when (flag_long='1') else '0';
	dataBufferOut( 574) <= dataBufferIn(2546) when (flag_long='1') else '0';
	dataBufferOut( 575) <= dataBufferIn(3289) when (flag_long='1') else '0';
	dataBufferOut( 576) <= dataBufferIn(4032) when (flag_long='1') else '0';
	dataBufferOut( 577) <= dataBufferIn(4775) when (flag_long='1') else '0';
	dataBufferOut( 578) <= dataBufferIn(5518) when (flag_long='1') else '0';
	dataBufferOut( 579) <= dataBufferIn( 117) when (flag_long='1') else '0';
	dataBufferOut( 580) <= dataBufferIn( 860) when (flag_long='1') else '0';
	dataBufferOut( 581) <= dataBufferIn(1603) when (flag_long='1') else '0';
	dataBufferOut( 582) <= dataBufferIn(2346) when (flag_long='1') else '0';
	dataBufferOut( 583) <= dataBufferIn(3089) when (flag_long='1') else '0';
	dataBufferOut( 584) <= dataBufferIn(3832) when (flag_long='1') else '0';
	dataBufferOut( 585) <= dataBufferIn(4575) when (flag_long='1') else '0';
	dataBufferOut( 586) <= dataBufferIn(5318) when (flag_long='1') else '0';
	dataBufferOut( 587) <= dataBufferIn(6061) when (flag_long='1') else '0';
	dataBufferOut( 588) <= dataBufferIn( 660) when (flag_long='1') else '0';
	dataBufferOut( 589) <= dataBufferIn(1403) when (flag_long='1') else '0';
	dataBufferOut( 590) <= dataBufferIn(2146) when (flag_long='1') else '0';
	dataBufferOut( 591) <= dataBufferIn(2889) when (flag_long='1') else '0';
	dataBufferOut( 592) <= dataBufferIn(3632) when (flag_long='1') else '0';
	dataBufferOut( 593) <= dataBufferIn(4375) when (flag_long='1') else '0';
	dataBufferOut( 594) <= dataBufferIn(5118) when (flag_long='1') else '0';
	dataBufferOut( 595) <= dataBufferIn(5861) when (flag_long='1') else '0';
	dataBufferOut( 596) <= dataBufferIn( 460) when (flag_long='1') else '0';
	dataBufferOut( 597) <= dataBufferIn(1203) when (flag_long='1') else '0';
	dataBufferOut( 598) <= dataBufferIn(1946) when (flag_long='1') else '0';
	dataBufferOut( 599) <= dataBufferIn(2689) when (flag_long='1') else '0';
	dataBufferOut( 600) <= dataBufferIn(3432) when (flag_long='1') else '0';
	dataBufferOut( 601) <= dataBufferIn(4175) when (flag_long='1') else '0';
	dataBufferOut( 602) <= dataBufferIn(4918) when (flag_long='1') else '0';
	dataBufferOut( 603) <= dataBufferIn(5661) when (flag_long='1') else '0';
	dataBufferOut( 604) <= dataBufferIn( 260) when (flag_long='1') else '0';
	dataBufferOut( 605) <= dataBufferIn(1003) when (flag_long='1') else '0';
	dataBufferOut( 606) <= dataBufferIn(1746) when (flag_long='1') else '0';
	dataBufferOut( 607) <= dataBufferIn(2489) when (flag_long='1') else '0';
	dataBufferOut( 608) <= dataBufferIn(3232) when (flag_long='1') else '0';
	dataBufferOut( 609) <= dataBufferIn(3975) when (flag_long='1') else '0';
	dataBufferOut( 610) <= dataBufferIn(4718) when (flag_long='1') else '0';
	dataBufferOut( 611) <= dataBufferIn(5461) when (flag_long='1') else '0';
	dataBufferOut( 612) <= dataBufferIn(  60) when (flag_long='1') else '0';
	dataBufferOut( 613) <= dataBufferIn( 803) when (flag_long='1') else '0';
	dataBufferOut( 614) <= dataBufferIn(1546) when (flag_long='1') else '0';
	dataBufferOut( 615) <= dataBufferIn(2289) when (flag_long='1') else '0';
	dataBufferOut( 616) <= dataBufferIn(3032) when (flag_long='1') else '0';
	dataBufferOut( 617) <= dataBufferIn(3775) when (flag_long='1') else '0';
	dataBufferOut( 618) <= dataBufferIn(4518) when (flag_long='1') else '0';
	dataBufferOut( 619) <= dataBufferIn(5261) when (flag_long='1') else '0';
	dataBufferOut( 620) <= dataBufferIn(6004) when (flag_long='1') else '0';
	dataBufferOut( 621) <= dataBufferIn( 603) when (flag_long='1') else '0';
	dataBufferOut( 622) <= dataBufferIn(1346) when (flag_long='1') else '0';
	dataBufferOut( 623) <= dataBufferIn(2089) when (flag_long='1') else '0';
	dataBufferOut( 624) <= dataBufferIn(2832) when (flag_long='1') else '0';
	dataBufferOut( 625) <= dataBufferIn(3575) when (flag_long='1') else '0';
	dataBufferOut( 626) <= dataBufferIn(4318) when (flag_long='1') else '0';
	dataBufferOut( 627) <= dataBufferIn(5061) when (flag_long='1') else '0';
	dataBufferOut( 628) <= dataBufferIn(5804) when (flag_long='1') else '0';
	dataBufferOut( 629) <= dataBufferIn( 403) when (flag_long='1') else '0';
	dataBufferOut( 630) <= dataBufferIn(1146) when (flag_long='1') else '0';
	dataBufferOut( 631) <= dataBufferIn(1889) when (flag_long='1') else '0';
	dataBufferOut( 632) <= dataBufferIn(2632) when (flag_long='1') else '0';
	dataBufferOut( 633) <= dataBufferIn(3375) when (flag_long='1') else '0';
	dataBufferOut( 634) <= dataBufferIn(4118) when (flag_long='1') else '0';
	dataBufferOut( 635) <= dataBufferIn(4861) when (flag_long='1') else '0';
	dataBufferOut( 636) <= dataBufferIn(5604) when (flag_long='1') else '0';
	dataBufferOut( 637) <= dataBufferIn( 203) when (flag_long='1') else '0';
	dataBufferOut( 638) <= dataBufferIn( 946) when (flag_long='1') else '0';
	dataBufferOut( 639) <= dataBufferIn(1689) when (flag_long='1') else '0';
	dataBufferOut( 640) <= dataBufferIn(2432) when (flag_long='1') else '0';
	dataBufferOut( 641) <= dataBufferIn(3175) when (flag_long='1') else '0';
	dataBufferOut( 642) <= dataBufferIn(3918) when (flag_long='1') else '0';
	dataBufferOut( 643) <= dataBufferIn(4661) when (flag_long='1') else '0';
	dataBufferOut( 644) <= dataBufferIn(5404) when (flag_long='1') else '0';
	dataBufferOut( 645) <= dataBufferIn(   3) when (flag_long='1') else '0';
	dataBufferOut( 646) <= dataBufferIn( 746) when (flag_long='1') else '0';
	dataBufferOut( 647) <= dataBufferIn(1489) when (flag_long='1') else '0';
	dataBufferOut( 648) <= dataBufferIn(2232) when (flag_long='1') else '0';
	dataBufferOut( 649) <= dataBufferIn(2975) when (flag_long='1') else '0';
	dataBufferOut( 650) <= dataBufferIn(3718) when (flag_long='1') else '0';
	dataBufferOut( 651) <= dataBufferIn(4461) when (flag_long='1') else '0';
	dataBufferOut( 652) <= dataBufferIn(5204) when (flag_long='1') else '0';
	dataBufferOut( 653) <= dataBufferIn(5947) when (flag_long='1') else '0';
	dataBufferOut( 654) <= dataBufferIn( 546) when (flag_long='1') else '0';
	dataBufferOut( 655) <= dataBufferIn(1289) when (flag_long='1') else '0';
	dataBufferOut( 656) <= dataBufferIn(2032) when (flag_long='1') else '0';
	dataBufferOut( 657) <= dataBufferIn(2775) when (flag_long='1') else '0';
	dataBufferOut( 658) <= dataBufferIn(3518) when (flag_long='1') else '0';
	dataBufferOut( 659) <= dataBufferIn(4261) when (flag_long='1') else '0';
	dataBufferOut( 660) <= dataBufferIn(5004) when (flag_long='1') else '0';
	dataBufferOut( 661) <= dataBufferIn(5747) when (flag_long='1') else '0';
	dataBufferOut( 662) <= dataBufferIn( 346) when (flag_long='1') else '0';
	dataBufferOut( 663) <= dataBufferIn(1089) when (flag_long='1') else '0';
	dataBufferOut( 664) <= dataBufferIn(1832) when (flag_long='1') else '0';
	dataBufferOut( 665) <= dataBufferIn(2575) when (flag_long='1') else '0';
	dataBufferOut( 666) <= dataBufferIn(3318) when (flag_long='1') else '0';
	dataBufferOut( 667) <= dataBufferIn(4061) when (flag_long='1') else '0';
	dataBufferOut( 668) <= dataBufferIn(4804) when (flag_long='1') else '0';
	dataBufferOut( 669) <= dataBufferIn(5547) when (flag_long='1') else '0';
	dataBufferOut( 670) <= dataBufferIn( 146) when (flag_long='1') else '0';
	dataBufferOut( 671) <= dataBufferIn( 889) when (flag_long='1') else '0';
	dataBufferOut( 672) <= dataBufferIn(1632) when (flag_long='1') else '0';
	dataBufferOut( 673) <= dataBufferIn(2375) when (flag_long='1') else '0';
	dataBufferOut( 674) <= dataBufferIn(3118) when (flag_long='1') else '0';
	dataBufferOut( 675) <= dataBufferIn(3861) when (flag_long='1') else '0';
	dataBufferOut( 676) <= dataBufferIn(4604) when (flag_long='1') else '0';
	dataBufferOut( 677) <= dataBufferIn(5347) when (flag_long='1') else '0';
	dataBufferOut( 678) <= dataBufferIn(6090) when (flag_long='1') else '0';
	dataBufferOut( 679) <= dataBufferIn( 689) when (flag_long='1') else '0';
	dataBufferOut( 680) <= dataBufferIn(1432) when (flag_long='1') else '0';
	dataBufferOut( 681) <= dataBufferIn(2175) when (flag_long='1') else '0';
	dataBufferOut( 682) <= dataBufferIn(2918) when (flag_long='1') else '0';
	dataBufferOut( 683) <= dataBufferIn(3661) when (flag_long='1') else '0';
	dataBufferOut( 684) <= dataBufferIn(4404) when (flag_long='1') else '0';
	dataBufferOut( 685) <= dataBufferIn(5147) when (flag_long='1') else '0';
	dataBufferOut( 686) <= dataBufferIn(5890) when (flag_long='1') else '0';
	dataBufferOut( 687) <= dataBufferIn( 489) when (flag_long='1') else '0';
	dataBufferOut( 688) <= dataBufferIn(1232) when (flag_long='1') else '0';
	dataBufferOut( 689) <= dataBufferIn(1975) when (flag_long='1') else '0';
	dataBufferOut( 690) <= dataBufferIn(2718) when (flag_long='1') else '0';
	dataBufferOut( 691) <= dataBufferIn(3461) when (flag_long='1') else '0';
	dataBufferOut( 692) <= dataBufferIn(4204) when (flag_long='1') else '0';
	dataBufferOut( 693) <= dataBufferIn(4947) when (flag_long='1') else '0';
	dataBufferOut( 694) <= dataBufferIn(5690) when (flag_long='1') else '0';
	dataBufferOut( 695) <= dataBufferIn( 289) when (flag_long='1') else '0';
	dataBufferOut( 696) <= dataBufferIn(1032) when (flag_long='1') else '0';
	dataBufferOut( 697) <= dataBufferIn(1775) when (flag_long='1') else '0';
	dataBufferOut( 698) <= dataBufferIn(2518) when (flag_long='1') else '0';
	dataBufferOut( 699) <= dataBufferIn(3261) when (flag_long='1') else '0';
	dataBufferOut( 700) <= dataBufferIn(4004) when (flag_long='1') else '0';
	dataBufferOut( 701) <= dataBufferIn(4747) when (flag_long='1') else '0';
	dataBufferOut( 702) <= dataBufferIn(5490) when (flag_long='1') else '0';
	dataBufferOut( 703) <= dataBufferIn(  89) when (flag_long='1') else '0';
	dataBufferOut( 704) <= dataBufferIn( 832) when (flag_long='1') else '0';
	dataBufferOut( 705) <= dataBufferIn(1575) when (flag_long='1') else '0';
	dataBufferOut( 706) <= dataBufferIn(2318) when (flag_long='1') else '0';
	dataBufferOut( 707) <= dataBufferIn(3061) when (flag_long='1') else '0';
	dataBufferOut( 708) <= dataBufferIn(3804) when (flag_long='1') else '0';
	dataBufferOut( 709) <= dataBufferIn(4547) when (flag_long='1') else '0';
	dataBufferOut( 710) <= dataBufferIn(5290) when (flag_long='1') else '0';
	dataBufferOut( 711) <= dataBufferIn(6033) when (flag_long='1') else '0';
	dataBufferOut( 712) <= dataBufferIn( 632) when (flag_long='1') else '0';
	dataBufferOut( 713) <= dataBufferIn(1375) when (flag_long='1') else '0';
	dataBufferOut( 714) <= dataBufferIn(2118) when (flag_long='1') else '0';
	dataBufferOut( 715) <= dataBufferIn(2861) when (flag_long='1') else '0';
	dataBufferOut( 716) <= dataBufferIn(3604) when (flag_long='1') else '0';
	dataBufferOut( 717) <= dataBufferIn(4347) when (flag_long='1') else '0';
	dataBufferOut( 718) <= dataBufferIn(5090) when (flag_long='1') else '0';
	dataBufferOut( 719) <= dataBufferIn(5833) when (flag_long='1') else '0';
	dataBufferOut( 720) <= dataBufferIn( 432) when (flag_long='1') else '0';
	dataBufferOut( 721) <= dataBufferIn(1175) when (flag_long='1') else '0';
	dataBufferOut( 722) <= dataBufferIn(1918) when (flag_long='1') else '0';
	dataBufferOut( 723) <= dataBufferIn(2661) when (flag_long='1') else '0';
	dataBufferOut( 724) <= dataBufferIn(3404) when (flag_long='1') else '0';
	dataBufferOut( 725) <= dataBufferIn(4147) when (flag_long='1') else '0';
	dataBufferOut( 726) <= dataBufferIn(4890) when (flag_long='1') else '0';
	dataBufferOut( 727) <= dataBufferIn(5633) when (flag_long='1') else '0';
	dataBufferOut( 728) <= dataBufferIn( 232) when (flag_long='1') else '0';
	dataBufferOut( 729) <= dataBufferIn( 975) when (flag_long='1') else '0';
	dataBufferOut( 730) <= dataBufferIn(1718) when (flag_long='1') else '0';
	dataBufferOut( 731) <= dataBufferIn(2461) when (flag_long='1') else '0';
	dataBufferOut( 732) <= dataBufferIn(3204) when (flag_long='1') else '0';
	dataBufferOut( 733) <= dataBufferIn(3947) when (flag_long='1') else '0';
	dataBufferOut( 734) <= dataBufferIn(4690) when (flag_long='1') else '0';
	dataBufferOut( 735) <= dataBufferIn(5433) when (flag_long='1') else '0';
	dataBufferOut( 736) <= dataBufferIn(  32) when (flag_long='1') else '0';
	dataBufferOut( 737) <= dataBufferIn( 775) when (flag_long='1') else '0';
	dataBufferOut( 738) <= dataBufferIn(1518) when (flag_long='1') else '0';
	dataBufferOut( 739) <= dataBufferIn(2261) when (flag_long='1') else '0';
	dataBufferOut( 740) <= dataBufferIn(3004) when (flag_long='1') else '0';
	dataBufferOut( 741) <= dataBufferIn(3747) when (flag_long='1') else '0';
	dataBufferOut( 742) <= dataBufferIn(4490) when (flag_long='1') else '0';
	dataBufferOut( 743) <= dataBufferIn(5233) when (flag_long='1') else '0';
	dataBufferOut( 744) <= dataBufferIn(5976) when (flag_long='1') else '0';
	dataBufferOut( 745) <= dataBufferIn( 575) when (flag_long='1') else '0';
	dataBufferOut( 746) <= dataBufferIn(1318) when (flag_long='1') else '0';
	dataBufferOut( 747) <= dataBufferIn(2061) when (flag_long='1') else '0';
	dataBufferOut( 748) <= dataBufferIn(2804) when (flag_long='1') else '0';
	dataBufferOut( 749) <= dataBufferIn(3547) when (flag_long='1') else '0';
	dataBufferOut( 750) <= dataBufferIn(4290) when (flag_long='1') else '0';
	dataBufferOut( 751) <= dataBufferIn(5033) when (flag_long='1') else '0';
	dataBufferOut( 752) <= dataBufferIn(5776) when (flag_long='1') else '0';
	dataBufferOut( 753) <= dataBufferIn( 375) when (flag_long='1') else '0';
	dataBufferOut( 754) <= dataBufferIn(1118) when (flag_long='1') else '0';
	dataBufferOut( 755) <= dataBufferIn(1861) when (flag_long='1') else '0';
	dataBufferOut( 756) <= dataBufferIn(2604) when (flag_long='1') else '0';
	dataBufferOut( 757) <= dataBufferIn(3347) when (flag_long='1') else '0';
	dataBufferOut( 758) <= dataBufferIn(4090) when (flag_long='1') else '0';
	dataBufferOut( 759) <= dataBufferIn(4833) when (flag_long='1') else '0';
	dataBufferOut( 760) <= dataBufferIn(5576) when (flag_long='1') else '0';
	dataBufferOut( 761) <= dataBufferIn( 175) when (flag_long='1') else '0';
	dataBufferOut( 762) <= dataBufferIn( 918) when (flag_long='1') else '0';
	dataBufferOut( 763) <= dataBufferIn(1661) when (flag_long='1') else '0';
	dataBufferOut( 764) <= dataBufferIn(2404) when (flag_long='1') else '0';
	dataBufferOut( 765) <= dataBufferIn(3147) when (flag_long='1') else '0';
	dataBufferOut( 766) <= dataBufferIn(3890) when (flag_long='1') else '0';
	dataBufferOut( 767) <= dataBufferIn(4633) when (flag_long='1') else '0';
	dataBufferOut( 768) <= dataBufferIn(5376) when (flag_long='1') else '0';
	dataBufferOut( 769) <= dataBufferIn(6119) when (flag_long='1') else '0';
	dataBufferOut( 770) <= dataBufferIn( 718) when (flag_long='1') else '0';
	dataBufferOut( 771) <= dataBufferIn(1461) when (flag_long='1') else '0';
	dataBufferOut( 772) <= dataBufferIn(2204) when (flag_long='1') else '0';
	dataBufferOut( 773) <= dataBufferIn(2947) when (flag_long='1') else '0';
	dataBufferOut( 774) <= dataBufferIn(3690) when (flag_long='1') else '0';
	dataBufferOut( 775) <= dataBufferIn(4433) when (flag_long='1') else '0';
	dataBufferOut( 776) <= dataBufferIn(5176) when (flag_long='1') else '0';
	dataBufferOut( 777) <= dataBufferIn(5919) when (flag_long='1') else '0';
	dataBufferOut( 778) <= dataBufferIn( 518) when (flag_long='1') else '0';
	dataBufferOut( 779) <= dataBufferIn(1261) when (flag_long='1') else '0';
	dataBufferOut( 780) <= dataBufferIn(2004) when (flag_long='1') else '0';
	dataBufferOut( 781) <= dataBufferIn(2747) when (flag_long='1') else '0';
	dataBufferOut( 782) <= dataBufferIn(3490) when (flag_long='1') else '0';
	dataBufferOut( 783) <= dataBufferIn(4233) when (flag_long='1') else '0';
	dataBufferOut( 784) <= dataBufferIn(4976) when (flag_long='1') else '0';
	dataBufferOut( 785) <= dataBufferIn(5719) when (flag_long='1') else '0';
	dataBufferOut( 786) <= dataBufferIn( 318) when (flag_long='1') else '0';
	dataBufferOut( 787) <= dataBufferIn(1061) when (flag_long='1') else '0';
	dataBufferOut( 788) <= dataBufferIn(1804) when (flag_long='1') else '0';
	dataBufferOut( 789) <= dataBufferIn(2547) when (flag_long='1') else '0';
	dataBufferOut( 790) <= dataBufferIn(3290) when (flag_long='1') else '0';
	dataBufferOut( 791) <= dataBufferIn(4033) when (flag_long='1') else '0';
	dataBufferOut( 792) <= dataBufferIn(4776) when (flag_long='1') else '0';
	dataBufferOut( 793) <= dataBufferIn(5519) when (flag_long='1') else '0';
	dataBufferOut( 794) <= dataBufferIn( 118) when (flag_long='1') else '0';
	dataBufferOut( 795) <= dataBufferIn( 861) when (flag_long='1') else '0';
	dataBufferOut( 796) <= dataBufferIn(1604) when (flag_long='1') else '0';
	dataBufferOut( 797) <= dataBufferIn(2347) when (flag_long='1') else '0';
	dataBufferOut( 798) <= dataBufferIn(3090) when (flag_long='1') else '0';
	dataBufferOut( 799) <= dataBufferIn(3833) when (flag_long='1') else '0';
	dataBufferOut( 800) <= dataBufferIn(4576) when (flag_long='1') else '0';
	dataBufferOut( 801) <= dataBufferIn(5319) when (flag_long='1') else '0';
	dataBufferOut( 802) <= dataBufferIn(6062) when (flag_long='1') else '0';
	dataBufferOut( 803) <= dataBufferIn( 661) when (flag_long='1') else '0';
	dataBufferOut( 804) <= dataBufferIn(1404) when (flag_long='1') else '0';
	dataBufferOut( 805) <= dataBufferIn(2147) when (flag_long='1') else '0';
	dataBufferOut( 806) <= dataBufferIn(2890) when (flag_long='1') else '0';
	dataBufferOut( 807) <= dataBufferIn(3633) when (flag_long='1') else '0';
	dataBufferOut( 808) <= dataBufferIn(4376) when (flag_long='1') else '0';
	dataBufferOut( 809) <= dataBufferIn(5119) when (flag_long='1') else '0';
	dataBufferOut( 810) <= dataBufferIn(5862) when (flag_long='1') else '0';
	dataBufferOut( 811) <= dataBufferIn( 461) when (flag_long='1') else '0';
	dataBufferOut( 812) <= dataBufferIn(1204) when (flag_long='1') else '0';
	dataBufferOut( 813) <= dataBufferIn(1947) when (flag_long='1') else '0';
	dataBufferOut( 814) <= dataBufferIn(2690) when (flag_long='1') else '0';
	dataBufferOut( 815) <= dataBufferIn(3433) when (flag_long='1') else '0';
	dataBufferOut( 816) <= dataBufferIn(4176) when (flag_long='1') else '0';
	dataBufferOut( 817) <= dataBufferIn(4919) when (flag_long='1') else '0';
	dataBufferOut( 818) <= dataBufferIn(5662) when (flag_long='1') else '0';
	dataBufferOut( 819) <= dataBufferIn( 261) when (flag_long='1') else '0';
	dataBufferOut( 820) <= dataBufferIn(1004) when (flag_long='1') else '0';
	dataBufferOut( 821) <= dataBufferIn(1747) when (flag_long='1') else '0';
	dataBufferOut( 822) <= dataBufferIn(2490) when (flag_long='1') else '0';
	dataBufferOut( 823) <= dataBufferIn(3233) when (flag_long='1') else '0';
	dataBufferOut( 824) <= dataBufferIn(3976) when (flag_long='1') else '0';
	dataBufferOut( 825) <= dataBufferIn(4719) when (flag_long='1') else '0';
	dataBufferOut( 826) <= dataBufferIn(5462) when (flag_long='1') else '0';
	dataBufferOut( 827) <= dataBufferIn(  61) when (flag_long='1') else '0';
	dataBufferOut( 828) <= dataBufferIn( 804) when (flag_long='1') else '0';
	dataBufferOut( 829) <= dataBufferIn(1547) when (flag_long='1') else '0';
	dataBufferOut( 830) <= dataBufferIn(2290) when (flag_long='1') else '0';
	dataBufferOut( 831) <= dataBufferIn(3033) when (flag_long='1') else '0';
	dataBufferOut( 832) <= dataBufferIn(3776) when (flag_long='1') else '0';
	dataBufferOut( 833) <= dataBufferIn(4519) when (flag_long='1') else '0';
	dataBufferOut( 834) <= dataBufferIn(5262) when (flag_long='1') else '0';
	dataBufferOut( 835) <= dataBufferIn(6005) when (flag_long='1') else '0';
	dataBufferOut( 836) <= dataBufferIn( 604) when (flag_long='1') else '0';
	dataBufferOut( 837) <= dataBufferIn(1347) when (flag_long='1') else '0';
	dataBufferOut( 838) <= dataBufferIn(2090) when (flag_long='1') else '0';
	dataBufferOut( 839) <= dataBufferIn(2833) when (flag_long='1') else '0';
	dataBufferOut( 840) <= dataBufferIn(3576) when (flag_long='1') else '0';
	dataBufferOut( 841) <= dataBufferIn(4319) when (flag_long='1') else '0';
	dataBufferOut( 842) <= dataBufferIn(5062) when (flag_long='1') else '0';
	dataBufferOut( 843) <= dataBufferIn(5805) when (flag_long='1') else '0';
	dataBufferOut( 844) <= dataBufferIn( 404) when (flag_long='1') else '0';
	dataBufferOut( 845) <= dataBufferIn(1147) when (flag_long='1') else '0';
	dataBufferOut( 846) <= dataBufferIn(1890) when (flag_long='1') else '0';
	dataBufferOut( 847) <= dataBufferIn(2633) when (flag_long='1') else '0';
	dataBufferOut( 848) <= dataBufferIn(3376) when (flag_long='1') else '0';
	dataBufferOut( 849) <= dataBufferIn(4119) when (flag_long='1') else '0';
	dataBufferOut( 850) <= dataBufferIn(4862) when (flag_long='1') else '0';
	dataBufferOut( 851) <= dataBufferIn(5605) when (flag_long='1') else '0';
	dataBufferOut( 852) <= dataBufferIn( 204) when (flag_long='1') else '0';
	dataBufferOut( 853) <= dataBufferIn( 947) when (flag_long='1') else '0';
	dataBufferOut( 854) <= dataBufferIn(1690) when (flag_long='1') else '0';
	dataBufferOut( 855) <= dataBufferIn(2433) when (flag_long='1') else '0';
	dataBufferOut( 856) <= dataBufferIn(3176) when (flag_long='1') else '0';
	dataBufferOut( 857) <= dataBufferIn(3919) when (flag_long='1') else '0';
	dataBufferOut( 858) <= dataBufferIn(4662) when (flag_long='1') else '0';
	dataBufferOut( 859) <= dataBufferIn(5405) when (flag_long='1') else '0';
	dataBufferOut( 860) <= dataBufferIn(   4) when (flag_long='1') else '0';
	dataBufferOut( 861) <= dataBufferIn( 747) when (flag_long='1') else '0';
	dataBufferOut( 862) <= dataBufferIn(1490) when (flag_long='1') else '0';
	dataBufferOut( 863) <= dataBufferIn(2233) when (flag_long='1') else '0';
	dataBufferOut( 864) <= dataBufferIn(2976) when (flag_long='1') else '0';
	dataBufferOut( 865) <= dataBufferIn(3719) when (flag_long='1') else '0';
	dataBufferOut( 866) <= dataBufferIn(4462) when (flag_long='1') else '0';
	dataBufferOut( 867) <= dataBufferIn(5205) when (flag_long='1') else '0';
	dataBufferOut( 868) <= dataBufferIn(5948) when (flag_long='1') else '0';
	dataBufferOut( 869) <= dataBufferIn( 547) when (flag_long='1') else '0';
	dataBufferOut( 870) <= dataBufferIn(1290) when (flag_long='1') else '0';
	dataBufferOut( 871) <= dataBufferIn(2033) when (flag_long='1') else '0';
	dataBufferOut( 872) <= dataBufferIn(2776) when (flag_long='1') else '0';
	dataBufferOut( 873) <= dataBufferIn(3519) when (flag_long='1') else '0';
	dataBufferOut( 874) <= dataBufferIn(4262) when (flag_long='1') else '0';
	dataBufferOut( 875) <= dataBufferIn(5005) when (flag_long='1') else '0';
	dataBufferOut( 876) <= dataBufferIn(5748) when (flag_long='1') else '0';
	dataBufferOut( 877) <= dataBufferIn( 347) when (flag_long='1') else '0';
	dataBufferOut( 878) <= dataBufferIn(1090) when (flag_long='1') else '0';
	dataBufferOut( 879) <= dataBufferIn(1833) when (flag_long='1') else '0';
	dataBufferOut( 880) <= dataBufferIn(2576) when (flag_long='1') else '0';
	dataBufferOut( 881) <= dataBufferIn(3319) when (flag_long='1') else '0';
	dataBufferOut( 882) <= dataBufferIn(4062) when (flag_long='1') else '0';
	dataBufferOut( 883) <= dataBufferIn(4805) when (flag_long='1') else '0';
	dataBufferOut( 884) <= dataBufferIn(5548) when (flag_long='1') else '0';
	dataBufferOut( 885) <= dataBufferIn( 147) when (flag_long='1') else '0';
	dataBufferOut( 886) <= dataBufferIn( 890) when (flag_long='1') else '0';
	dataBufferOut( 887) <= dataBufferIn(1633) when (flag_long='1') else '0';
	dataBufferOut( 888) <= dataBufferIn(2376) when (flag_long='1') else '0';
	dataBufferOut( 889) <= dataBufferIn(3119) when (flag_long='1') else '0';
	dataBufferOut( 890) <= dataBufferIn(3862) when (flag_long='1') else '0';
	dataBufferOut( 891) <= dataBufferIn(4605) when (flag_long='1') else '0';
	dataBufferOut( 892) <= dataBufferIn(5348) when (flag_long='1') else '0';
	dataBufferOut( 893) <= dataBufferIn(6091) when (flag_long='1') else '0';
	dataBufferOut( 894) <= dataBufferIn( 690) when (flag_long='1') else '0';
	dataBufferOut( 895) <= dataBufferIn(1433) when (flag_long='1') else '0';
	dataBufferOut( 896) <= dataBufferIn(2176) when (flag_long='1') else '0';
	dataBufferOut( 897) <= dataBufferIn(2919) when (flag_long='1') else '0';
	dataBufferOut( 898) <= dataBufferIn(3662) when (flag_long='1') else '0';
	dataBufferOut( 899) <= dataBufferIn(4405) when (flag_long='1') else '0';
	dataBufferOut( 900) <= dataBufferIn(5148) when (flag_long='1') else '0';
	dataBufferOut( 901) <= dataBufferIn(5891) when (flag_long='1') else '0';
	dataBufferOut( 902) <= dataBufferIn( 490) when (flag_long='1') else '0';
	dataBufferOut( 903) <= dataBufferIn(1233) when (flag_long='1') else '0';
	dataBufferOut( 904) <= dataBufferIn(1976) when (flag_long='1') else '0';
	dataBufferOut( 905) <= dataBufferIn(2719) when (flag_long='1') else '0';
	dataBufferOut( 906) <= dataBufferIn(3462) when (flag_long='1') else '0';
	dataBufferOut( 907) <= dataBufferIn(4205) when (flag_long='1') else '0';
	dataBufferOut( 908) <= dataBufferIn(4948) when (flag_long='1') else '0';
	dataBufferOut( 909) <= dataBufferIn(5691) when (flag_long='1') else '0';
	dataBufferOut( 910) <= dataBufferIn( 290) when (flag_long='1') else '0';
	dataBufferOut( 911) <= dataBufferIn(1033) when (flag_long='1') else '0';
	dataBufferOut( 912) <= dataBufferIn(1776) when (flag_long='1') else '0';
	dataBufferOut( 913) <= dataBufferIn(2519) when (flag_long='1') else '0';
	dataBufferOut( 914) <= dataBufferIn(3262) when (flag_long='1') else '0';
	dataBufferOut( 915) <= dataBufferIn(4005) when (flag_long='1') else '0';
	dataBufferOut( 916) <= dataBufferIn(4748) when (flag_long='1') else '0';
	dataBufferOut( 917) <= dataBufferIn(5491) when (flag_long='1') else '0';
	dataBufferOut( 918) <= dataBufferIn(  90) when (flag_long='1') else '0';
	dataBufferOut( 919) <= dataBufferIn( 833) when (flag_long='1') else '0';
	dataBufferOut( 920) <= dataBufferIn(1576) when (flag_long='1') else '0';
	dataBufferOut( 921) <= dataBufferIn(2319) when (flag_long='1') else '0';
	dataBufferOut( 922) <= dataBufferIn(3062) when (flag_long='1') else '0';
	dataBufferOut( 923) <= dataBufferIn(3805) when (flag_long='1') else '0';
	dataBufferOut( 924) <= dataBufferIn(4548) when (flag_long='1') else '0';
	dataBufferOut( 925) <= dataBufferIn(5291) when (flag_long='1') else '0';
	dataBufferOut( 926) <= dataBufferIn(6034) when (flag_long='1') else '0';
	dataBufferOut( 927) <= dataBufferIn( 633) when (flag_long='1') else '0';
	dataBufferOut( 928) <= dataBufferIn(1376) when (flag_long='1') else '0';
	dataBufferOut( 929) <= dataBufferIn(2119) when (flag_long='1') else '0';
	dataBufferOut( 930) <= dataBufferIn(2862) when (flag_long='1') else '0';
	dataBufferOut( 931) <= dataBufferIn(3605) when (flag_long='1') else '0';
	dataBufferOut( 932) <= dataBufferIn(4348) when (flag_long='1') else '0';
	dataBufferOut( 933) <= dataBufferIn(5091) when (flag_long='1') else '0';
	dataBufferOut( 934) <= dataBufferIn(5834) when (flag_long='1') else '0';
	dataBufferOut( 935) <= dataBufferIn( 433) when (flag_long='1') else '0';
	dataBufferOut( 936) <= dataBufferIn(1176) when (flag_long='1') else '0';
	dataBufferOut( 937) <= dataBufferIn(1919) when (flag_long='1') else '0';
	dataBufferOut( 938) <= dataBufferIn(2662) when (flag_long='1') else '0';
	dataBufferOut( 939) <= dataBufferIn(3405) when (flag_long='1') else '0';
	dataBufferOut( 940) <= dataBufferIn(4148) when (flag_long='1') else '0';
	dataBufferOut( 941) <= dataBufferIn(4891) when (flag_long='1') else '0';
	dataBufferOut( 942) <= dataBufferIn(5634) when (flag_long='1') else '0';
	dataBufferOut( 943) <= dataBufferIn( 233) when (flag_long='1') else '0';
	dataBufferOut( 944) <= dataBufferIn( 976) when (flag_long='1') else '0';
	dataBufferOut( 945) <= dataBufferIn(1719) when (flag_long='1') else '0';
	dataBufferOut( 946) <= dataBufferIn(2462) when (flag_long='1') else '0';
	dataBufferOut( 947) <= dataBufferIn(3205) when (flag_long='1') else '0';
	dataBufferOut( 948) <= dataBufferIn(3948) when (flag_long='1') else '0';
	dataBufferOut( 949) <= dataBufferIn(4691) when (flag_long='1') else '0';
	dataBufferOut( 950) <= dataBufferIn(5434) when (flag_long='1') else '0';
	dataBufferOut( 951) <= dataBufferIn(  33) when (flag_long='1') else '0';
	dataBufferOut( 952) <= dataBufferIn( 776) when (flag_long='1') else '0';
	dataBufferOut( 953) <= dataBufferIn(1519) when (flag_long='1') else '0';
	dataBufferOut( 954) <= dataBufferIn(2262) when (flag_long='1') else '0';
	dataBufferOut( 955) <= dataBufferIn(3005) when (flag_long='1') else '0';
	dataBufferOut( 956) <= dataBufferIn(3748) when (flag_long='1') else '0';
	dataBufferOut( 957) <= dataBufferIn(4491) when (flag_long='1') else '0';
	dataBufferOut( 958) <= dataBufferIn(5234) when (flag_long='1') else '0';
	dataBufferOut( 959) <= dataBufferIn(5977) when (flag_long='1') else '0';
	dataBufferOut( 960) <= dataBufferIn( 576) when (flag_long='1') else '0';
	dataBufferOut( 961) <= dataBufferIn(1319) when (flag_long='1') else '0';
	dataBufferOut( 962) <= dataBufferIn(2062) when (flag_long='1') else '0';
	dataBufferOut( 963) <= dataBufferIn(2805) when (flag_long='1') else '0';
	dataBufferOut( 964) <= dataBufferIn(3548) when (flag_long='1') else '0';
	dataBufferOut( 965) <= dataBufferIn(4291) when (flag_long='1') else '0';
	dataBufferOut( 966) <= dataBufferIn(5034) when (flag_long='1') else '0';
	dataBufferOut( 967) <= dataBufferIn(5777) when (flag_long='1') else '0';
	dataBufferOut( 968) <= dataBufferIn( 376) when (flag_long='1') else '0';
	dataBufferOut( 969) <= dataBufferIn(1119) when (flag_long='1') else '0';
	dataBufferOut( 970) <= dataBufferIn(1862) when (flag_long='1') else '0';
	dataBufferOut( 971) <= dataBufferIn(2605) when (flag_long='1') else '0';
	dataBufferOut( 972) <= dataBufferIn(3348) when (flag_long='1') else '0';
	dataBufferOut( 973) <= dataBufferIn(4091) when (flag_long='1') else '0';
	dataBufferOut( 974) <= dataBufferIn(4834) when (flag_long='1') else '0';
	dataBufferOut( 975) <= dataBufferIn(5577) when (flag_long='1') else '0';
	dataBufferOut( 976) <= dataBufferIn( 176) when (flag_long='1') else '0';
	dataBufferOut( 977) <= dataBufferIn( 919) when (flag_long='1') else '0';
	dataBufferOut( 978) <= dataBufferIn(1662) when (flag_long='1') else '0';
	dataBufferOut( 979) <= dataBufferIn(2405) when (flag_long='1') else '0';
	dataBufferOut( 980) <= dataBufferIn(3148) when (flag_long='1') else '0';
	dataBufferOut( 981) <= dataBufferIn(3891) when (flag_long='1') else '0';
	dataBufferOut( 982) <= dataBufferIn(4634) when (flag_long='1') else '0';
	dataBufferOut( 983) <= dataBufferIn(5377) when (flag_long='1') else '0';
	dataBufferOut( 984) <= dataBufferIn(6120) when (flag_long='1') else '0';
	dataBufferOut( 985) <= dataBufferIn( 719) when (flag_long='1') else '0';
	dataBufferOut( 986) <= dataBufferIn(1462) when (flag_long='1') else '0';
	dataBufferOut( 987) <= dataBufferIn(2205) when (flag_long='1') else '0';
	dataBufferOut( 988) <= dataBufferIn(2948) when (flag_long='1') else '0';
	dataBufferOut( 989) <= dataBufferIn(3691) when (flag_long='1') else '0';
	dataBufferOut( 990) <= dataBufferIn(4434) when (flag_long='1') else '0';
	dataBufferOut( 991) <= dataBufferIn(5177) when (flag_long='1') else '0';
	dataBufferOut( 992) <= dataBufferIn(5920) when (flag_long='1') else '0';
	dataBufferOut( 993) <= dataBufferIn( 519) when (flag_long='1') else '0';
	dataBufferOut( 994) <= dataBufferIn(1262) when (flag_long='1') else '0';
	dataBufferOut( 995) <= dataBufferIn(2005) when (flag_long='1') else '0';
	dataBufferOut( 996) <= dataBufferIn(2748) when (flag_long='1') else '0';
	dataBufferOut( 997) <= dataBufferIn(3491) when (flag_long='1') else '0';
	dataBufferOut( 998) <= dataBufferIn(4234) when (flag_long='1') else '0';
	dataBufferOut( 999) <= dataBufferIn(4977) when (flag_long='1') else '0';
	dataBufferOut(1000) <= dataBufferIn(5720) when (flag_long='1') else '0';
	dataBufferOut(1001) <= dataBufferIn( 319) when (flag_long='1') else '0';
	dataBufferOut(1002) <= dataBufferIn(1062) when (flag_long='1') else '0';
	dataBufferOut(1003) <= dataBufferIn(1805) when (flag_long='1') else '0';
	dataBufferOut(1004) <= dataBufferIn(2548) when (flag_long='1') else '0';
	dataBufferOut(1005) <= dataBufferIn(3291) when (flag_long='1') else '0';
	dataBufferOut(1006) <= dataBufferIn(4034) when (flag_long='1') else '0';
	dataBufferOut(1007) <= dataBufferIn(4777) when (flag_long='1') else '0';
	dataBufferOut(1008) <= dataBufferIn(5520) when (flag_long='1') else '0';
	dataBufferOut(1009) <= dataBufferIn( 119) when (flag_long='1') else '0';
	dataBufferOut(1010) <= dataBufferIn( 862) when (flag_long='1') else '0';
	dataBufferOut(1011) <= dataBufferIn(1605) when (flag_long='1') else '0';
	dataBufferOut(1012) <= dataBufferIn(2348) when (flag_long='1') else '0';
	dataBufferOut(1013) <= dataBufferIn(3091) when (flag_long='1') else '0';
	dataBufferOut(1014) <= dataBufferIn(3834) when (flag_long='1') else '0';
	dataBufferOut(1015) <= dataBufferIn(4577) when (flag_long='1') else '0';
	dataBufferOut(1016) <= dataBufferIn(5320) when (flag_long='1') else '0';
	dataBufferOut(1017) <= dataBufferIn(6063) when (flag_long='1') else '0';
	dataBufferOut(1018) <= dataBufferIn( 662) when (flag_long='1') else '0';
	dataBufferOut(1019) <= dataBufferIn(1405) when (flag_long='1') else '0';
	dataBufferOut(1020) <= dataBufferIn(2148) when (flag_long='1') else '0';
	dataBufferOut(1021) <= dataBufferIn(2891) when (flag_long='1') else '0';
	dataBufferOut(1022) <= dataBufferIn(3634) when (flag_long='1') else '0';
	dataBufferOut(1023) <= dataBufferIn(4377) when (flag_long='1') else '0';
	dataBufferOut(1024) <= dataBufferIn(5120) when (flag_long='1') else '0';
	dataBufferOut(1025) <= dataBufferIn(5863) when (flag_long='1') else '0';
	dataBufferOut(1026) <= dataBufferIn( 462) when (flag_long='1') else '0';
	dataBufferOut(1027) <= dataBufferIn(1205) when (flag_long='1') else '0';
	dataBufferOut(1028) <= dataBufferIn(1948) when (flag_long='1') else '0';
	dataBufferOut(1029) <= dataBufferIn(2691) when (flag_long='1') else '0';
	dataBufferOut(1030) <= dataBufferIn(3434) when (flag_long='1') else '0';
	dataBufferOut(1031) <= dataBufferIn(4177) when (flag_long='1') else '0';
	dataBufferOut(1032) <= dataBufferIn(4920) when (flag_long='1') else '0';
	dataBufferOut(1033) <= dataBufferIn(5663) when (flag_long='1') else '0';
	dataBufferOut(1034) <= dataBufferIn( 262) when (flag_long='1') else '0';
	dataBufferOut(1035) <= dataBufferIn(1005) when (flag_long='1') else '0';
	dataBufferOut(1036) <= dataBufferIn(1748) when (flag_long='1') else '0';
	dataBufferOut(1037) <= dataBufferIn(2491) when (flag_long='1') else '0';
	dataBufferOut(1038) <= dataBufferIn(3234) when (flag_long='1') else '0';
	dataBufferOut(1039) <= dataBufferIn(3977) when (flag_long='1') else '0';
	dataBufferOut(1040) <= dataBufferIn(4720) when (flag_long='1') else '0';
	dataBufferOut(1041) <= dataBufferIn(5463) when (flag_long='1') else '0';
	dataBufferOut(1042) <= dataBufferIn(  62) when (flag_long='1') else '0';
	dataBufferOut(1043) <= dataBufferIn( 805) when (flag_long='1') else '0';
	dataBufferOut(1044) <= dataBufferIn(1548) when (flag_long='1') else '0';
	dataBufferOut(1045) <= dataBufferIn(2291) when (flag_long='1') else '0';
	dataBufferOut(1046) <= dataBufferIn(3034) when (flag_long='1') else '0';
	dataBufferOut(1047) <= dataBufferIn(3777) when (flag_long='1') else '0';
	dataBufferOut(1048) <= dataBufferIn(4520) when (flag_long='1') else '0';
	dataBufferOut(1049) <= dataBufferIn(5263) when (flag_long='1') else '0';
	dataBufferOut(1050) <= dataBufferIn(6006) when (flag_long='1') else '0';
	dataBufferOut(1051) <= dataBufferIn( 605) when (flag_long='1') else '0';
	dataBufferOut(1052) <= dataBufferIn(1348) when (flag_long='1') else '0';
	dataBufferOut(1053) <= dataBufferIn(2091) when (flag_long='1') else '0';
	dataBufferOut(1054) <= dataBufferIn(2834) when (flag_long='1') else '0';
	dataBufferOut(1055) <= dataBufferIn(3577) when (flag_long='1') else '0';
	dataBufferOut(1056) <= dataBufferIn(4320) when (flag_long='1') else '0';
	dataBufferOut(1057) <= dataBufferIn(5063) when (flag_long='1') else '0';
	dataBufferOut(1058) <= dataBufferIn(5806) when (flag_long='1') else '0';
	dataBufferOut(1059) <= dataBufferIn( 405) when (flag_long='1') else '0';
	dataBufferOut(1060) <= dataBufferIn(1148) when (flag_long='1') else '0';
	dataBufferOut(1061) <= dataBufferIn(1891) when (flag_long='1') else '0';
	dataBufferOut(1062) <= dataBufferIn(2634) when (flag_long='1') else '0';
	dataBufferOut(1063) <= dataBufferIn(3377) when (flag_long='1') else '0';
	dataBufferOut(1064) <= dataBufferIn(4120) when (flag_long='1') else '0';
	dataBufferOut(1065) <= dataBufferIn(4863) when (flag_long='1') else '0';
	dataBufferOut(1066) <= dataBufferIn(5606) when (flag_long='1') else '0';
	dataBufferOut(1067) <= dataBufferIn( 205) when (flag_long='1') else '0';
	dataBufferOut(1068) <= dataBufferIn( 948) when (flag_long='1') else '0';
	dataBufferOut(1069) <= dataBufferIn(1691) when (flag_long='1') else '0';
	dataBufferOut(1070) <= dataBufferIn(2434) when (flag_long='1') else '0';
	dataBufferOut(1071) <= dataBufferIn(3177) when (flag_long='1') else '0';
	dataBufferOut(1072) <= dataBufferIn(3920) when (flag_long='1') else '0';
	dataBufferOut(1073) <= dataBufferIn(4663) when (flag_long='1') else '0';
	dataBufferOut(1074) <= dataBufferIn(5406) when (flag_long='1') else '0';
	dataBufferOut(1075) <= dataBufferIn(   5) when (flag_long='1') else '0';
	dataBufferOut(1076) <= dataBufferIn( 748) when (flag_long='1') else '0';
	dataBufferOut(1077) <= dataBufferIn(1491) when (flag_long='1') else '0';
	dataBufferOut(1078) <= dataBufferIn(2234) when (flag_long='1') else '0';
	dataBufferOut(1079) <= dataBufferIn(2977) when (flag_long='1') else '0';
	dataBufferOut(1080) <= dataBufferIn(3720) when (flag_long='1') else '0';
	dataBufferOut(1081) <= dataBufferIn(4463) when (flag_long='1') else '0';
	dataBufferOut(1082) <= dataBufferIn(5206) when (flag_long='1') else '0';
	dataBufferOut(1083) <= dataBufferIn(5949) when (flag_long='1') else '0';
	dataBufferOut(1084) <= dataBufferIn( 548) when (flag_long='1') else '0';
	dataBufferOut(1085) <= dataBufferIn(1291) when (flag_long='1') else '0';
	dataBufferOut(1086) <= dataBufferIn(2034) when (flag_long='1') else '0';
	dataBufferOut(1087) <= dataBufferIn(2777) when (flag_long='1') else '0';
	dataBufferOut(1088) <= dataBufferIn(3520) when (flag_long='1') else '0';
	dataBufferOut(1089) <= dataBufferIn(4263) when (flag_long='1') else '0';
	dataBufferOut(1090) <= dataBufferIn(5006) when (flag_long='1') else '0';
	dataBufferOut(1091) <= dataBufferIn(5749) when (flag_long='1') else '0';
	dataBufferOut(1092) <= dataBufferIn( 348) when (flag_long='1') else '0';
	dataBufferOut(1093) <= dataBufferIn(1091) when (flag_long='1') else '0';
	dataBufferOut(1094) <= dataBufferIn(1834) when (flag_long='1') else '0';
	dataBufferOut(1095) <= dataBufferIn(2577) when (flag_long='1') else '0';
	dataBufferOut(1096) <= dataBufferIn(3320) when (flag_long='1') else '0';
	dataBufferOut(1097) <= dataBufferIn(4063) when (flag_long='1') else '0';
	dataBufferOut(1098) <= dataBufferIn(4806) when (flag_long='1') else '0';
	dataBufferOut(1099) <= dataBufferIn(5549) when (flag_long='1') else '0';
	dataBufferOut(1100) <= dataBufferIn( 148) when (flag_long='1') else '0';
	dataBufferOut(1101) <= dataBufferIn( 891) when (flag_long='1') else '0';
	dataBufferOut(1102) <= dataBufferIn(1634) when (flag_long='1') else '0';
	dataBufferOut(1103) <= dataBufferIn(2377) when (flag_long='1') else '0';
	dataBufferOut(1104) <= dataBufferIn(3120) when (flag_long='1') else '0';
	dataBufferOut(1105) <= dataBufferIn(3863) when (flag_long='1') else '0';
	dataBufferOut(1106) <= dataBufferIn(4606) when (flag_long='1') else '0';
	dataBufferOut(1107) <= dataBufferIn(5349) when (flag_long='1') else '0';
	dataBufferOut(1108) <= dataBufferIn(6092) when (flag_long='1') else '0';
	dataBufferOut(1109) <= dataBufferIn( 691) when (flag_long='1') else '0';
	dataBufferOut(1110) <= dataBufferIn(1434) when (flag_long='1') else '0';
	dataBufferOut(1111) <= dataBufferIn(2177) when (flag_long='1') else '0';
	dataBufferOut(1112) <= dataBufferIn(2920) when (flag_long='1') else '0';
	dataBufferOut(1113) <= dataBufferIn(3663) when (flag_long='1') else '0';
	dataBufferOut(1114) <= dataBufferIn(4406) when (flag_long='1') else '0';
	dataBufferOut(1115) <= dataBufferIn(5149) when (flag_long='1') else '0';
	dataBufferOut(1116) <= dataBufferIn(5892) when (flag_long='1') else '0';
	dataBufferOut(1117) <= dataBufferIn( 491) when (flag_long='1') else '0';
	dataBufferOut(1118) <= dataBufferIn(1234) when (flag_long='1') else '0';
	dataBufferOut(1119) <= dataBufferIn(1977) when (flag_long='1') else '0';
	dataBufferOut(1120) <= dataBufferIn(2720) when (flag_long='1') else '0';
	dataBufferOut(1121) <= dataBufferIn(3463) when (flag_long='1') else '0';
	dataBufferOut(1122) <= dataBufferIn(4206) when (flag_long='1') else '0';
	dataBufferOut(1123) <= dataBufferIn(4949) when (flag_long='1') else '0';
	dataBufferOut(1124) <= dataBufferIn(5692) when (flag_long='1') else '0';
	dataBufferOut(1125) <= dataBufferIn( 291) when (flag_long='1') else '0';
	dataBufferOut(1126) <= dataBufferIn(1034) when (flag_long='1') else '0';
	dataBufferOut(1127) <= dataBufferIn(1777) when (flag_long='1') else '0';
	dataBufferOut(1128) <= dataBufferIn(2520) when (flag_long='1') else '0';
	dataBufferOut(1129) <= dataBufferIn(3263) when (flag_long='1') else '0';
	dataBufferOut(1130) <= dataBufferIn(4006) when (flag_long='1') else '0';
	dataBufferOut(1131) <= dataBufferIn(4749) when (flag_long='1') else '0';
	dataBufferOut(1132) <= dataBufferIn(5492) when (flag_long='1') else '0';
	dataBufferOut(1133) <= dataBufferIn(  91) when (flag_long='1') else '0';
	dataBufferOut(1134) <= dataBufferIn( 834) when (flag_long='1') else '0';
	dataBufferOut(1135) <= dataBufferIn(1577) when (flag_long='1') else '0';
	dataBufferOut(1136) <= dataBufferIn(2320) when (flag_long='1') else '0';
	dataBufferOut(1137) <= dataBufferIn(3063) when (flag_long='1') else '0';
	dataBufferOut(1138) <= dataBufferIn(3806) when (flag_long='1') else '0';
	dataBufferOut(1139) <= dataBufferIn(4549) when (flag_long='1') else '0';
	dataBufferOut(1140) <= dataBufferIn(5292) when (flag_long='1') else '0';
	dataBufferOut(1141) <= dataBufferIn(6035) when (flag_long='1') else '0';
	dataBufferOut(1142) <= dataBufferIn( 634) when (flag_long='1') else '0';
	dataBufferOut(1143) <= dataBufferIn(1377) when (flag_long='1') else '0';
	dataBufferOut(1144) <= dataBufferIn(2120) when (flag_long='1') else '0';
	dataBufferOut(1145) <= dataBufferIn(2863) when (flag_long='1') else '0';
	dataBufferOut(1146) <= dataBufferIn(3606) when (flag_long='1') else '0';
	dataBufferOut(1147) <= dataBufferIn(4349) when (flag_long='1') else '0';
	dataBufferOut(1148) <= dataBufferIn(5092) when (flag_long='1') else '0';
	dataBufferOut(1149) <= dataBufferIn(5835) when (flag_long='1') else '0';
	dataBufferOut(1150) <= dataBufferIn( 434) when (flag_long='1') else '0';
	dataBufferOut(1151) <= dataBufferIn(1177) when (flag_long='1') else '0';
	dataBufferOut(1152) <= dataBufferIn(1920) when (flag_long='1') else '0';
	dataBufferOut(1153) <= dataBufferIn(2663) when (flag_long='1') else '0';
	dataBufferOut(1154) <= dataBufferIn(3406) when (flag_long='1') else '0';
	dataBufferOut(1155) <= dataBufferIn(4149) when (flag_long='1') else '0';
	dataBufferOut(1156) <= dataBufferIn(4892) when (flag_long='1') else '0';
	dataBufferOut(1157) <= dataBufferIn(5635) when (flag_long='1') else '0';
	dataBufferOut(1158) <= dataBufferIn( 234) when (flag_long='1') else '0';
	dataBufferOut(1159) <= dataBufferIn( 977) when (flag_long='1') else '0';
	dataBufferOut(1160) <= dataBufferIn(1720) when (flag_long='1') else '0';
	dataBufferOut(1161) <= dataBufferIn(2463) when (flag_long='1') else '0';
	dataBufferOut(1162) <= dataBufferIn(3206) when (flag_long='1') else '0';
	dataBufferOut(1163) <= dataBufferIn(3949) when (flag_long='1') else '0';
	dataBufferOut(1164) <= dataBufferIn(4692) when (flag_long='1') else '0';
	dataBufferOut(1165) <= dataBufferIn(5435) when (flag_long='1') else '0';
	dataBufferOut(1166) <= dataBufferIn(  34) when (flag_long='1') else '0';
	dataBufferOut(1167) <= dataBufferIn( 777) when (flag_long='1') else '0';
	dataBufferOut(1168) <= dataBufferIn(1520) when (flag_long='1') else '0';
	dataBufferOut(1169) <= dataBufferIn(2263) when (flag_long='1') else '0';
	dataBufferOut(1170) <= dataBufferIn(3006) when (flag_long='1') else '0';
	dataBufferOut(1171) <= dataBufferIn(3749) when (flag_long='1') else '0';
	dataBufferOut(1172) <= dataBufferIn(4492) when (flag_long='1') else '0';
	dataBufferOut(1173) <= dataBufferIn(5235) when (flag_long='1') else '0';
	dataBufferOut(1174) <= dataBufferIn(5978) when (flag_long='1') else '0';
	dataBufferOut(1175) <= dataBufferIn( 577) when (flag_long='1') else '0';
	dataBufferOut(1176) <= dataBufferIn(1320) when (flag_long='1') else '0';
	dataBufferOut(1177) <= dataBufferIn(2063) when (flag_long='1') else '0';
	dataBufferOut(1178) <= dataBufferIn(2806) when (flag_long='1') else '0';
	dataBufferOut(1179) <= dataBufferIn(3549) when (flag_long='1') else '0';
	dataBufferOut(1180) <= dataBufferIn(4292) when (flag_long='1') else '0';
	dataBufferOut(1181) <= dataBufferIn(5035) when (flag_long='1') else '0';
	dataBufferOut(1182) <= dataBufferIn(5778) when (flag_long='1') else '0';
	dataBufferOut(1183) <= dataBufferIn( 377) when (flag_long='1') else '0';
	dataBufferOut(1184) <= dataBufferIn(1120) when (flag_long='1') else '0';
	dataBufferOut(1185) <= dataBufferIn(1863) when (flag_long='1') else '0';
	dataBufferOut(1186) <= dataBufferIn(2606) when (flag_long='1') else '0';
	dataBufferOut(1187) <= dataBufferIn(3349) when (flag_long='1') else '0';
	dataBufferOut(1188) <= dataBufferIn(4092) when (flag_long='1') else '0';
	dataBufferOut(1189) <= dataBufferIn(4835) when (flag_long='1') else '0';
	dataBufferOut(1190) <= dataBufferIn(5578) when (flag_long='1') else '0';
	dataBufferOut(1191) <= dataBufferIn( 177) when (flag_long='1') else '0';
	dataBufferOut(1192) <= dataBufferIn( 920) when (flag_long='1') else '0';
	dataBufferOut(1193) <= dataBufferIn(1663) when (flag_long='1') else '0';
	dataBufferOut(1194) <= dataBufferIn(2406) when (flag_long='1') else '0';
	dataBufferOut(1195) <= dataBufferIn(3149) when (flag_long='1') else '0';
	dataBufferOut(1196) <= dataBufferIn(3892) when (flag_long='1') else '0';
	dataBufferOut(1197) <= dataBufferIn(4635) when (flag_long='1') else '0';
	dataBufferOut(1198) <= dataBufferIn(5378) when (flag_long='1') else '0';
	dataBufferOut(1199) <= dataBufferIn(6121) when (flag_long='1') else '0';
	dataBufferOut(1200) <= dataBufferIn( 720) when (flag_long='1') else '0';
	dataBufferOut(1201) <= dataBufferIn(1463) when (flag_long='1') else '0';
	dataBufferOut(1202) <= dataBufferIn(2206) when (flag_long='1') else '0';
	dataBufferOut(1203) <= dataBufferIn(2949) when (flag_long='1') else '0';
	dataBufferOut(1204) <= dataBufferIn(3692) when (flag_long='1') else '0';
	dataBufferOut(1205) <= dataBufferIn(4435) when (flag_long='1') else '0';
	dataBufferOut(1206) <= dataBufferIn(5178) when (flag_long='1') else '0';
	dataBufferOut(1207) <= dataBufferIn(5921) when (flag_long='1') else '0';
	dataBufferOut(1208) <= dataBufferIn( 520) when (flag_long='1') else '0';
	dataBufferOut(1209) <= dataBufferIn(1263) when (flag_long='1') else '0';
	dataBufferOut(1210) <= dataBufferIn(2006) when (flag_long='1') else '0';
	dataBufferOut(1211) <= dataBufferIn(2749) when (flag_long='1') else '0';
	dataBufferOut(1212) <= dataBufferIn(3492) when (flag_long='1') else '0';
	dataBufferOut(1213) <= dataBufferIn(4235) when (flag_long='1') else '0';
	dataBufferOut(1214) <= dataBufferIn(4978) when (flag_long='1') else '0';
	dataBufferOut(1215) <= dataBufferIn(5721) when (flag_long='1') else '0';
	dataBufferOut(1216) <= dataBufferIn( 320) when (flag_long='1') else '0';
	dataBufferOut(1217) <= dataBufferIn(1063) when (flag_long='1') else '0';
	dataBufferOut(1218) <= dataBufferIn(1806) when (flag_long='1') else '0';
	dataBufferOut(1219) <= dataBufferIn(2549) when (flag_long='1') else '0';
	dataBufferOut(1220) <= dataBufferIn(3292) when (flag_long='1') else '0';
	dataBufferOut(1221) <= dataBufferIn(4035) when (flag_long='1') else '0';
	dataBufferOut(1222) <= dataBufferIn(4778) when (flag_long='1') else '0';
	dataBufferOut(1223) <= dataBufferIn(5521) when (flag_long='1') else '0';
	dataBufferOut(1224) <= dataBufferIn( 120) when (flag_long='1') else '0';
	dataBufferOut(1225) <= dataBufferIn( 863) when (flag_long='1') else '0';
	dataBufferOut(1226) <= dataBufferIn(1606) when (flag_long='1') else '0';
	dataBufferOut(1227) <= dataBufferIn(2349) when (flag_long='1') else '0';
	dataBufferOut(1228) <= dataBufferIn(3092) when (flag_long='1') else '0';
	dataBufferOut(1229) <= dataBufferIn(3835) when (flag_long='1') else '0';
	dataBufferOut(1230) <= dataBufferIn(4578) when (flag_long='1') else '0';
	dataBufferOut(1231) <= dataBufferIn(5321) when (flag_long='1') else '0';
	dataBufferOut(1232) <= dataBufferIn(6064) when (flag_long='1') else '0';
	dataBufferOut(1233) <= dataBufferIn( 663) when (flag_long='1') else '0';
	dataBufferOut(1234) <= dataBufferIn(1406) when (flag_long='1') else '0';
	dataBufferOut(1235) <= dataBufferIn(2149) when (flag_long='1') else '0';
	dataBufferOut(1236) <= dataBufferIn(2892) when (flag_long='1') else '0';
	dataBufferOut(1237) <= dataBufferIn(3635) when (flag_long='1') else '0';
	dataBufferOut(1238) <= dataBufferIn(4378) when (flag_long='1') else '0';
	dataBufferOut(1239) <= dataBufferIn(5121) when (flag_long='1') else '0';
	dataBufferOut(1240) <= dataBufferIn(5864) when (flag_long='1') else '0';
	dataBufferOut(1241) <= dataBufferIn( 463) when (flag_long='1') else '0';
	dataBufferOut(1242) <= dataBufferIn(1206) when (flag_long='1') else '0';
	dataBufferOut(1243) <= dataBufferIn(1949) when (flag_long='1') else '0';
	dataBufferOut(1244) <= dataBufferIn(2692) when (flag_long='1') else '0';
	dataBufferOut(1245) <= dataBufferIn(3435) when (flag_long='1') else '0';
	dataBufferOut(1246) <= dataBufferIn(4178) when (flag_long='1') else '0';
	dataBufferOut(1247) <= dataBufferIn(4921) when (flag_long='1') else '0';
	dataBufferOut(1248) <= dataBufferIn(5664) when (flag_long='1') else '0';
	dataBufferOut(1249) <= dataBufferIn( 263) when (flag_long='1') else '0';
	dataBufferOut(1250) <= dataBufferIn(1006) when (flag_long='1') else '0';
	dataBufferOut(1251) <= dataBufferIn(1749) when (flag_long='1') else '0';
	dataBufferOut(1252) <= dataBufferIn(2492) when (flag_long='1') else '0';
	dataBufferOut(1253) <= dataBufferIn(3235) when (flag_long='1') else '0';
	dataBufferOut(1254) <= dataBufferIn(3978) when (flag_long='1') else '0';
	dataBufferOut(1255) <= dataBufferIn(4721) when (flag_long='1') else '0';
	dataBufferOut(1256) <= dataBufferIn(5464) when (flag_long='1') else '0';
	dataBufferOut(1257) <= dataBufferIn(  63) when (flag_long='1') else '0';
	dataBufferOut(1258) <= dataBufferIn( 806) when (flag_long='1') else '0';
	dataBufferOut(1259) <= dataBufferIn(1549) when (flag_long='1') else '0';
	dataBufferOut(1260) <= dataBufferIn(2292) when (flag_long='1') else '0';
	dataBufferOut(1261) <= dataBufferIn(3035) when (flag_long='1') else '0';
	dataBufferOut(1262) <= dataBufferIn(3778) when (flag_long='1') else '0';
	dataBufferOut(1263) <= dataBufferIn(4521) when (flag_long='1') else '0';
	dataBufferOut(1264) <= dataBufferIn(5264) when (flag_long='1') else '0';
	dataBufferOut(1265) <= dataBufferIn(6007) when (flag_long='1') else '0';
	dataBufferOut(1266) <= dataBufferIn( 606) when (flag_long='1') else '0';
	dataBufferOut(1267) <= dataBufferIn(1349) when (flag_long='1') else '0';
	dataBufferOut(1268) <= dataBufferIn(2092) when (flag_long='1') else '0';
	dataBufferOut(1269) <= dataBufferIn(2835) when (flag_long='1') else '0';
	dataBufferOut(1270) <= dataBufferIn(3578) when (flag_long='1') else '0';
	dataBufferOut(1271) <= dataBufferIn(4321) when (flag_long='1') else '0';
	dataBufferOut(1272) <= dataBufferIn(5064) when (flag_long='1') else '0';
	dataBufferOut(1273) <= dataBufferIn(5807) when (flag_long='1') else '0';
	dataBufferOut(1274) <= dataBufferIn( 406) when (flag_long='1') else '0';
	dataBufferOut(1275) <= dataBufferIn(1149) when (flag_long='1') else '0';
	dataBufferOut(1276) <= dataBufferIn(1892) when (flag_long='1') else '0';
	dataBufferOut(1277) <= dataBufferIn(2635) when (flag_long='1') else '0';
	dataBufferOut(1278) <= dataBufferIn(3378) when (flag_long='1') else '0';
	dataBufferOut(1279) <= dataBufferIn(4121) when (flag_long='1') else '0';
	dataBufferOut(1280) <= dataBufferIn(4864) when (flag_long='1') else '0';
	dataBufferOut(1281) <= dataBufferIn(5607) when (flag_long='1') else '0';
	dataBufferOut(1282) <= dataBufferIn( 206) when (flag_long='1') else '0';
	dataBufferOut(1283) <= dataBufferIn( 949) when (flag_long='1') else '0';
	dataBufferOut(1284) <= dataBufferIn(1692) when (flag_long='1') else '0';
	dataBufferOut(1285) <= dataBufferIn(2435) when (flag_long='1') else '0';
	dataBufferOut(1286) <= dataBufferIn(3178) when (flag_long='1') else '0';
	dataBufferOut(1287) <= dataBufferIn(3921) when (flag_long='1') else '0';
	dataBufferOut(1288) <= dataBufferIn(4664) when (flag_long='1') else '0';
	dataBufferOut(1289) <= dataBufferIn(5407) when (flag_long='1') else '0';
	dataBufferOut(1290) <= dataBufferIn(   6) when (flag_long='1') else '0';
	dataBufferOut(1291) <= dataBufferIn( 749) when (flag_long='1') else '0';
	dataBufferOut(1292) <= dataBufferIn(1492) when (flag_long='1') else '0';
	dataBufferOut(1293) <= dataBufferIn(2235) when (flag_long='1') else '0';
	dataBufferOut(1294) <= dataBufferIn(2978) when (flag_long='1') else '0';
	dataBufferOut(1295) <= dataBufferIn(3721) when (flag_long='1') else '0';
	dataBufferOut(1296) <= dataBufferIn(4464) when (flag_long='1') else '0';
	dataBufferOut(1297) <= dataBufferIn(5207) when (flag_long='1') else '0';
	dataBufferOut(1298) <= dataBufferIn(5950) when (flag_long='1') else '0';
	dataBufferOut(1299) <= dataBufferIn( 549) when (flag_long='1') else '0';
	dataBufferOut(1300) <= dataBufferIn(1292) when (flag_long='1') else '0';
	dataBufferOut(1301) <= dataBufferIn(2035) when (flag_long='1') else '0';
	dataBufferOut(1302) <= dataBufferIn(2778) when (flag_long='1') else '0';
	dataBufferOut(1303) <= dataBufferIn(3521) when (flag_long='1') else '0';
	dataBufferOut(1304) <= dataBufferIn(4264) when (flag_long='1') else '0';
	dataBufferOut(1305) <= dataBufferIn(5007) when (flag_long='1') else '0';
	dataBufferOut(1306) <= dataBufferIn(5750) when (flag_long='1') else '0';
	dataBufferOut(1307) <= dataBufferIn( 349) when (flag_long='1') else '0';
	dataBufferOut(1308) <= dataBufferIn(1092) when (flag_long='1') else '0';
	dataBufferOut(1309) <= dataBufferIn(1835) when (flag_long='1') else '0';
	dataBufferOut(1310) <= dataBufferIn(2578) when (flag_long='1') else '0';
	dataBufferOut(1311) <= dataBufferIn(3321) when (flag_long='1') else '0';
	dataBufferOut(1312) <= dataBufferIn(4064) when (flag_long='1') else '0';
	dataBufferOut(1313) <= dataBufferIn(4807) when (flag_long='1') else '0';
	dataBufferOut(1314) <= dataBufferIn(5550) when (flag_long='1') else '0';
	dataBufferOut(1315) <= dataBufferIn( 149) when (flag_long='1') else '0';
	dataBufferOut(1316) <= dataBufferIn( 892) when (flag_long='1') else '0';
	dataBufferOut(1317) <= dataBufferIn(1635) when (flag_long='1') else '0';
	dataBufferOut(1318) <= dataBufferIn(2378) when (flag_long='1') else '0';
	dataBufferOut(1319) <= dataBufferIn(3121) when (flag_long='1') else '0';
	dataBufferOut(1320) <= dataBufferIn(3864) when (flag_long='1') else '0';
	dataBufferOut(1321) <= dataBufferIn(4607) when (flag_long='1') else '0';
	dataBufferOut(1322) <= dataBufferIn(5350) when (flag_long='1') else '0';
	dataBufferOut(1323) <= dataBufferIn(6093) when (flag_long='1') else '0';
	dataBufferOut(1324) <= dataBufferIn( 692) when (flag_long='1') else '0';
	dataBufferOut(1325) <= dataBufferIn(1435) when (flag_long='1') else '0';
	dataBufferOut(1326) <= dataBufferIn(2178) when (flag_long='1') else '0';
	dataBufferOut(1327) <= dataBufferIn(2921) when (flag_long='1') else '0';
	dataBufferOut(1328) <= dataBufferIn(3664) when (flag_long='1') else '0';
	dataBufferOut(1329) <= dataBufferIn(4407) when (flag_long='1') else '0';
	dataBufferOut(1330) <= dataBufferIn(5150) when (flag_long='1') else '0';
	dataBufferOut(1331) <= dataBufferIn(5893) when (flag_long='1') else '0';
	dataBufferOut(1332) <= dataBufferIn( 492) when (flag_long='1') else '0';
	dataBufferOut(1333) <= dataBufferIn(1235) when (flag_long='1') else '0';
	dataBufferOut(1334) <= dataBufferIn(1978) when (flag_long='1') else '0';
	dataBufferOut(1335) <= dataBufferIn(2721) when (flag_long='1') else '0';
	dataBufferOut(1336) <= dataBufferIn(3464) when (flag_long='1') else '0';
	dataBufferOut(1337) <= dataBufferIn(4207) when (flag_long='1') else '0';
	dataBufferOut(1338) <= dataBufferIn(4950) when (flag_long='1') else '0';
	dataBufferOut(1339) <= dataBufferIn(5693) when (flag_long='1') else '0';
	dataBufferOut(1340) <= dataBufferIn( 292) when (flag_long='1') else '0';
	dataBufferOut(1341) <= dataBufferIn(1035) when (flag_long='1') else '0';
	dataBufferOut(1342) <= dataBufferIn(1778) when (flag_long='1') else '0';
	dataBufferOut(1343) <= dataBufferIn(2521) when (flag_long='1') else '0';
	dataBufferOut(1344) <= dataBufferIn(3264) when (flag_long='1') else '0';
	dataBufferOut(1345) <= dataBufferIn(4007) when (flag_long='1') else '0';
	dataBufferOut(1346) <= dataBufferIn(4750) when (flag_long='1') else '0';
	dataBufferOut(1347) <= dataBufferIn(5493) when (flag_long='1') else '0';
	dataBufferOut(1348) <= dataBufferIn(  92) when (flag_long='1') else '0';
	dataBufferOut(1349) <= dataBufferIn( 835) when (flag_long='1') else '0';
	dataBufferOut(1350) <= dataBufferIn(1578) when (flag_long='1') else '0';
	dataBufferOut(1351) <= dataBufferIn(2321) when (flag_long='1') else '0';
	dataBufferOut(1352) <= dataBufferIn(3064) when (flag_long='1') else '0';
	dataBufferOut(1353) <= dataBufferIn(3807) when (flag_long='1') else '0';
	dataBufferOut(1354) <= dataBufferIn(4550) when (flag_long='1') else '0';
	dataBufferOut(1355) <= dataBufferIn(5293) when (flag_long='1') else '0';
	dataBufferOut(1356) <= dataBufferIn(6036) when (flag_long='1') else '0';
	dataBufferOut(1357) <= dataBufferIn( 635) when (flag_long='1') else '0';
	dataBufferOut(1358) <= dataBufferIn(1378) when (flag_long='1') else '0';
	dataBufferOut(1359) <= dataBufferIn(2121) when (flag_long='1') else '0';
	dataBufferOut(1360) <= dataBufferIn(2864) when (flag_long='1') else '0';
	dataBufferOut(1361) <= dataBufferIn(3607) when (flag_long='1') else '0';
	dataBufferOut(1362) <= dataBufferIn(4350) when (flag_long='1') else '0';
	dataBufferOut(1363) <= dataBufferIn(5093) when (flag_long='1') else '0';
	dataBufferOut(1364) <= dataBufferIn(5836) when (flag_long='1') else '0';
	dataBufferOut(1365) <= dataBufferIn( 435) when (flag_long='1') else '0';
	dataBufferOut(1366) <= dataBufferIn(1178) when (flag_long='1') else '0';
	dataBufferOut(1367) <= dataBufferIn(1921) when (flag_long='1') else '0';
	dataBufferOut(1368) <= dataBufferIn(2664) when (flag_long='1') else '0';
	dataBufferOut(1369) <= dataBufferIn(3407) when (flag_long='1') else '0';
	dataBufferOut(1370) <= dataBufferIn(4150) when (flag_long='1') else '0';
	dataBufferOut(1371) <= dataBufferIn(4893) when (flag_long='1') else '0';
	dataBufferOut(1372) <= dataBufferIn(5636) when (flag_long='1') else '0';
	dataBufferOut(1373) <= dataBufferIn( 235) when (flag_long='1') else '0';
	dataBufferOut(1374) <= dataBufferIn( 978) when (flag_long='1') else '0';
	dataBufferOut(1375) <= dataBufferIn(1721) when (flag_long='1') else '0';
	dataBufferOut(1376) <= dataBufferIn(2464) when (flag_long='1') else '0';
	dataBufferOut(1377) <= dataBufferIn(3207) when (flag_long='1') else '0';
	dataBufferOut(1378) <= dataBufferIn(3950) when (flag_long='1') else '0';
	dataBufferOut(1379) <= dataBufferIn(4693) when (flag_long='1') else '0';
	dataBufferOut(1380) <= dataBufferIn(5436) when (flag_long='1') else '0';
	dataBufferOut(1381) <= dataBufferIn(  35) when (flag_long='1') else '0';
	dataBufferOut(1382) <= dataBufferIn( 778) when (flag_long='1') else '0';
	dataBufferOut(1383) <= dataBufferIn(1521) when (flag_long='1') else '0';
	dataBufferOut(1384) <= dataBufferIn(2264) when (flag_long='1') else '0';
	dataBufferOut(1385) <= dataBufferIn(3007) when (flag_long='1') else '0';
	dataBufferOut(1386) <= dataBufferIn(3750) when (flag_long='1') else '0';
	dataBufferOut(1387) <= dataBufferIn(4493) when (flag_long='1') else '0';
	dataBufferOut(1388) <= dataBufferIn(5236) when (flag_long='1') else '0';
	dataBufferOut(1389) <= dataBufferIn(5979) when (flag_long='1') else '0';
	dataBufferOut(1390) <= dataBufferIn( 578) when (flag_long='1') else '0';
	dataBufferOut(1391) <= dataBufferIn(1321) when (flag_long='1') else '0';
	dataBufferOut(1392) <= dataBufferIn(2064) when (flag_long='1') else '0';
	dataBufferOut(1393) <= dataBufferIn(2807) when (flag_long='1') else '0';
	dataBufferOut(1394) <= dataBufferIn(3550) when (flag_long='1') else '0';
	dataBufferOut(1395) <= dataBufferIn(4293) when (flag_long='1') else '0';
	dataBufferOut(1396) <= dataBufferIn(5036) when (flag_long='1') else '0';
	dataBufferOut(1397) <= dataBufferIn(5779) when (flag_long='1') else '0';
	dataBufferOut(1398) <= dataBufferIn( 378) when (flag_long='1') else '0';
	dataBufferOut(1399) <= dataBufferIn(1121) when (flag_long='1') else '0';
	dataBufferOut(1400) <= dataBufferIn(1864) when (flag_long='1') else '0';
	dataBufferOut(1401) <= dataBufferIn(2607) when (flag_long='1') else '0';
	dataBufferOut(1402) <= dataBufferIn(3350) when (flag_long='1') else '0';
	dataBufferOut(1403) <= dataBufferIn(4093) when (flag_long='1') else '0';
	dataBufferOut(1404) <= dataBufferIn(4836) when (flag_long='1') else '0';
	dataBufferOut(1405) <= dataBufferIn(5579) when (flag_long='1') else '0';
	dataBufferOut(1406) <= dataBufferIn( 178) when (flag_long='1') else '0';
	dataBufferOut(1407) <= dataBufferIn( 921) when (flag_long='1') else '0';
	dataBufferOut(1408) <= dataBufferIn(1664) when (flag_long='1') else '0';
	dataBufferOut(1409) <= dataBufferIn(2407) when (flag_long='1') else '0';
	dataBufferOut(1410) <= dataBufferIn(3150) when (flag_long='1') else '0';
	dataBufferOut(1411) <= dataBufferIn(3893) when (flag_long='1') else '0';
	dataBufferOut(1412) <= dataBufferIn(4636) when (flag_long='1') else '0';
	dataBufferOut(1413) <= dataBufferIn(5379) when (flag_long='1') else '0';
	dataBufferOut(1414) <= dataBufferIn(6122) when (flag_long='1') else '0';
	dataBufferOut(1415) <= dataBufferIn( 721) when (flag_long='1') else '0';
	dataBufferOut(1416) <= dataBufferIn(1464) when (flag_long='1') else '0';
	dataBufferOut(1417) <= dataBufferIn(2207) when (flag_long='1') else '0';
	dataBufferOut(1418) <= dataBufferIn(2950) when (flag_long='1') else '0';
	dataBufferOut(1419) <= dataBufferIn(3693) when (flag_long='1') else '0';
	dataBufferOut(1420) <= dataBufferIn(4436) when (flag_long='1') else '0';
	dataBufferOut(1421) <= dataBufferIn(5179) when (flag_long='1') else '0';
	dataBufferOut(1422) <= dataBufferIn(5922) when (flag_long='1') else '0';
	dataBufferOut(1423) <= dataBufferIn( 521) when (flag_long='1') else '0';
	dataBufferOut(1424) <= dataBufferIn(1264) when (flag_long='1') else '0';
	dataBufferOut(1425) <= dataBufferIn(2007) when (flag_long='1') else '0';
	dataBufferOut(1426) <= dataBufferIn(2750) when (flag_long='1') else '0';
	dataBufferOut(1427) <= dataBufferIn(3493) when (flag_long='1') else '0';
	dataBufferOut(1428) <= dataBufferIn(4236) when (flag_long='1') else '0';
	dataBufferOut(1429) <= dataBufferIn(4979) when (flag_long='1') else '0';
	dataBufferOut(1430) <= dataBufferIn(5722) when (flag_long='1') else '0';
	dataBufferOut(1431) <= dataBufferIn( 321) when (flag_long='1') else '0';
	dataBufferOut(1432) <= dataBufferIn(1064) when (flag_long='1') else '0';
	dataBufferOut(1433) <= dataBufferIn(1807) when (flag_long='1') else '0';
	dataBufferOut(1434) <= dataBufferIn(2550) when (flag_long='1') else '0';
	dataBufferOut(1435) <= dataBufferIn(3293) when (flag_long='1') else '0';
	dataBufferOut(1436) <= dataBufferIn(4036) when (flag_long='1') else '0';
	dataBufferOut(1437) <= dataBufferIn(4779) when (flag_long='1') else '0';
	dataBufferOut(1438) <= dataBufferIn(5522) when (flag_long='1') else '0';
	dataBufferOut(1439) <= dataBufferIn( 121) when (flag_long='1') else '0';
	dataBufferOut(1440) <= dataBufferIn( 864) when (flag_long='1') else '0';
	dataBufferOut(1441) <= dataBufferIn(1607) when (flag_long='1') else '0';
	dataBufferOut(1442) <= dataBufferIn(2350) when (flag_long='1') else '0';
	dataBufferOut(1443) <= dataBufferIn(3093) when (flag_long='1') else '0';
	dataBufferOut(1444) <= dataBufferIn(3836) when (flag_long='1') else '0';
	dataBufferOut(1445) <= dataBufferIn(4579) when (flag_long='1') else '0';
	dataBufferOut(1446) <= dataBufferIn(5322) when (flag_long='1') else '0';
	dataBufferOut(1447) <= dataBufferIn(6065) when (flag_long='1') else '0';
	dataBufferOut(1448) <= dataBufferIn( 664) when (flag_long='1') else '0';
	dataBufferOut(1449) <= dataBufferIn(1407) when (flag_long='1') else '0';
	dataBufferOut(1450) <= dataBufferIn(2150) when (flag_long='1') else '0';
	dataBufferOut(1451) <= dataBufferIn(2893) when (flag_long='1') else '0';
	dataBufferOut(1452) <= dataBufferIn(3636) when (flag_long='1') else '0';
	dataBufferOut(1453) <= dataBufferIn(4379) when (flag_long='1') else '0';
	dataBufferOut(1454) <= dataBufferIn(5122) when (flag_long='1') else '0';
	dataBufferOut(1455) <= dataBufferIn(5865) when (flag_long='1') else '0';
	dataBufferOut(1456) <= dataBufferIn( 464) when (flag_long='1') else '0';
	dataBufferOut(1457) <= dataBufferIn(1207) when (flag_long='1') else '0';
	dataBufferOut(1458) <= dataBufferIn(1950) when (flag_long='1') else '0';
	dataBufferOut(1459) <= dataBufferIn(2693) when (flag_long='1') else '0';
	dataBufferOut(1460) <= dataBufferIn(3436) when (flag_long='1') else '0';
	dataBufferOut(1461) <= dataBufferIn(4179) when (flag_long='1') else '0';
	dataBufferOut(1462) <= dataBufferIn(4922) when (flag_long='1') else '0';
	dataBufferOut(1463) <= dataBufferIn(5665) when (flag_long='1') else '0';
	dataBufferOut(1464) <= dataBufferIn( 264) when (flag_long='1') else '0';
	dataBufferOut(1465) <= dataBufferIn(1007) when (flag_long='1') else '0';
	dataBufferOut(1466) <= dataBufferIn(1750) when (flag_long='1') else '0';
	dataBufferOut(1467) <= dataBufferIn(2493) when (flag_long='1') else '0';
	dataBufferOut(1468) <= dataBufferIn(3236) when (flag_long='1') else '0';
	dataBufferOut(1469) <= dataBufferIn(3979) when (flag_long='1') else '0';
	dataBufferOut(1470) <= dataBufferIn(4722) when (flag_long='1') else '0';
	dataBufferOut(1471) <= dataBufferIn(5465) when (flag_long='1') else '0';
	dataBufferOut(1472) <= dataBufferIn(  64) when (flag_long='1') else '0';
	dataBufferOut(1473) <= dataBufferIn( 807) when (flag_long='1') else '0';
	dataBufferOut(1474) <= dataBufferIn(1550) when (flag_long='1') else '0';
	dataBufferOut(1475) <= dataBufferIn(2293) when (flag_long='1') else '0';
	dataBufferOut(1476) <= dataBufferIn(3036) when (flag_long='1') else '0';
	dataBufferOut(1477) <= dataBufferIn(3779) when (flag_long='1') else '0';
	dataBufferOut(1478) <= dataBufferIn(4522) when (flag_long='1') else '0';
	dataBufferOut(1479) <= dataBufferIn(5265) when (flag_long='1') else '0';
	dataBufferOut(1480) <= dataBufferIn(6008) when (flag_long='1') else '0';
	dataBufferOut(1481) <= dataBufferIn( 607) when (flag_long='1') else '0';
	dataBufferOut(1482) <= dataBufferIn(1350) when (flag_long='1') else '0';
	dataBufferOut(1483) <= dataBufferIn(2093) when (flag_long='1') else '0';
	dataBufferOut(1484) <= dataBufferIn(2836) when (flag_long='1') else '0';
	dataBufferOut(1485) <= dataBufferIn(3579) when (flag_long='1') else '0';
	dataBufferOut(1486) <= dataBufferIn(4322) when (flag_long='1') else '0';
	dataBufferOut(1487) <= dataBufferIn(5065) when (flag_long='1') else '0';
	dataBufferOut(1488) <= dataBufferIn(5808) when (flag_long='1') else '0';
	dataBufferOut(1489) <= dataBufferIn( 407) when (flag_long='1') else '0';
	dataBufferOut(1490) <= dataBufferIn(1150) when (flag_long='1') else '0';
	dataBufferOut(1491) <= dataBufferIn(1893) when (flag_long='1') else '0';
	dataBufferOut(1492) <= dataBufferIn(2636) when (flag_long='1') else '0';
	dataBufferOut(1493) <= dataBufferIn(3379) when (flag_long='1') else '0';
	dataBufferOut(1494) <= dataBufferIn(4122) when (flag_long='1') else '0';
	dataBufferOut(1495) <= dataBufferIn(4865) when (flag_long='1') else '0';
	dataBufferOut(1496) <= dataBufferIn(5608) when (flag_long='1') else '0';
	dataBufferOut(1497) <= dataBufferIn( 207) when (flag_long='1') else '0';
	dataBufferOut(1498) <= dataBufferIn( 950) when (flag_long='1') else '0';
	dataBufferOut(1499) <= dataBufferIn(1693) when (flag_long='1') else '0';
	dataBufferOut(1500) <= dataBufferIn(2436) when (flag_long='1') else '0';
	dataBufferOut(1501) <= dataBufferIn(3179) when (flag_long='1') else '0';
	dataBufferOut(1502) <= dataBufferIn(3922) when (flag_long='1') else '0';
	dataBufferOut(1503) <= dataBufferIn(4665) when (flag_long='1') else '0';
	dataBufferOut(1504) <= dataBufferIn(5408) when (flag_long='1') else '0';
	dataBufferOut(1505) <= dataBufferIn(   7) when (flag_long='1') else '0';
	dataBufferOut(1506) <= dataBufferIn( 750) when (flag_long='1') else '0';
	dataBufferOut(1507) <= dataBufferIn(1493) when (flag_long='1') else '0';
	dataBufferOut(1508) <= dataBufferIn(2236) when (flag_long='1') else '0';
	dataBufferOut(1509) <= dataBufferIn(2979) when (flag_long='1') else '0';
	dataBufferOut(1510) <= dataBufferIn(3722) when (flag_long='1') else '0';
	dataBufferOut(1511) <= dataBufferIn(4465) when (flag_long='1') else '0';
	dataBufferOut(1512) <= dataBufferIn(5208) when (flag_long='1') else '0';
	dataBufferOut(1513) <= dataBufferIn(5951) when (flag_long='1') else '0';
	dataBufferOut(1514) <= dataBufferIn( 550) when (flag_long='1') else '0';
	dataBufferOut(1515) <= dataBufferIn(1293) when (flag_long='1') else '0';
	dataBufferOut(1516) <= dataBufferIn(2036) when (flag_long='1') else '0';
	dataBufferOut(1517) <= dataBufferIn(2779) when (flag_long='1') else '0';
	dataBufferOut(1518) <= dataBufferIn(3522) when (flag_long='1') else '0';
	dataBufferOut(1519) <= dataBufferIn(4265) when (flag_long='1') else '0';
	dataBufferOut(1520) <= dataBufferIn(5008) when (flag_long='1') else '0';
	dataBufferOut(1521) <= dataBufferIn(5751) when (flag_long='1') else '0';
	dataBufferOut(1522) <= dataBufferIn( 350) when (flag_long='1') else '0';
	dataBufferOut(1523) <= dataBufferIn(1093) when (flag_long='1') else '0';
	dataBufferOut(1524) <= dataBufferIn(1836) when (flag_long='1') else '0';
	dataBufferOut(1525) <= dataBufferIn(2579) when (flag_long='1') else '0';
	dataBufferOut(1526) <= dataBufferIn(3322) when (flag_long='1') else '0';
	dataBufferOut(1527) <= dataBufferIn(4065) when (flag_long='1') else '0';
	dataBufferOut(1528) <= dataBufferIn(4808) when (flag_long='1') else '0';
	dataBufferOut(1529) <= dataBufferIn(5551) when (flag_long='1') else '0';
	dataBufferOut(1530) <= dataBufferIn( 150) when (flag_long='1') else '0';
	dataBufferOut(1531) <= dataBufferIn( 893) when (flag_long='1') else '0';
	dataBufferOut(1532) <= dataBufferIn(1636) when (flag_long='1') else '0';
	dataBufferOut(1533) <= dataBufferIn(2379) when (flag_long='1') else '0';
	dataBufferOut(1534) <= dataBufferIn(3122) when (flag_long='1') else '0';
	dataBufferOut(1535) <= dataBufferIn(3865) when (flag_long='1') else '0';
	dataBufferOut(1536) <= dataBufferIn(4608) when (flag_long='1') else '0';
	dataBufferOut(1537) <= dataBufferIn(5351) when (flag_long='1') else '0';
	dataBufferOut(1538) <= dataBufferIn(6094) when (flag_long='1') else '0';
	dataBufferOut(1539) <= dataBufferIn( 693) when (flag_long='1') else '0';
	dataBufferOut(1540) <= dataBufferIn(1436) when (flag_long='1') else '0';
	dataBufferOut(1541) <= dataBufferIn(2179) when (flag_long='1') else '0';
	dataBufferOut(1542) <= dataBufferIn(2922) when (flag_long='1') else '0';
	dataBufferOut(1543) <= dataBufferIn(3665) when (flag_long='1') else '0';
	dataBufferOut(1544) <= dataBufferIn(4408) when (flag_long='1') else '0';
	dataBufferOut(1545) <= dataBufferIn(5151) when (flag_long='1') else '0';
	dataBufferOut(1546) <= dataBufferIn(5894) when (flag_long='1') else '0';
	dataBufferOut(1547) <= dataBufferIn( 493) when (flag_long='1') else '0';
	dataBufferOut(1548) <= dataBufferIn(1236) when (flag_long='1') else '0';
	dataBufferOut(1549) <= dataBufferIn(1979) when (flag_long='1') else '0';
	dataBufferOut(1550) <= dataBufferIn(2722) when (flag_long='1') else '0';
	dataBufferOut(1551) <= dataBufferIn(3465) when (flag_long='1') else '0';
	dataBufferOut(1552) <= dataBufferIn(4208) when (flag_long='1') else '0';
	dataBufferOut(1553) <= dataBufferIn(4951) when (flag_long='1') else '0';
	dataBufferOut(1554) <= dataBufferIn(5694) when (flag_long='1') else '0';
	dataBufferOut(1555) <= dataBufferIn( 293) when (flag_long='1') else '0';
	dataBufferOut(1556) <= dataBufferIn(1036) when (flag_long='1') else '0';
	dataBufferOut(1557) <= dataBufferIn(1779) when (flag_long='1') else '0';
	dataBufferOut(1558) <= dataBufferIn(2522) when (flag_long='1') else '0';
	dataBufferOut(1559) <= dataBufferIn(3265) when (flag_long='1') else '0';
	dataBufferOut(1560) <= dataBufferIn(4008) when (flag_long='1') else '0';
	dataBufferOut(1561) <= dataBufferIn(4751) when (flag_long='1') else '0';
	dataBufferOut(1562) <= dataBufferIn(5494) when (flag_long='1') else '0';
	dataBufferOut(1563) <= dataBufferIn(  93) when (flag_long='1') else '0';
	dataBufferOut(1564) <= dataBufferIn( 836) when (flag_long='1') else '0';
	dataBufferOut(1565) <= dataBufferIn(1579) when (flag_long='1') else '0';
	dataBufferOut(1566) <= dataBufferIn(2322) when (flag_long='1') else '0';
	dataBufferOut(1567) <= dataBufferIn(3065) when (flag_long='1') else '0';
	dataBufferOut(1568) <= dataBufferIn(3808) when (flag_long='1') else '0';
	dataBufferOut(1569) <= dataBufferIn(4551) when (flag_long='1') else '0';
	dataBufferOut(1570) <= dataBufferIn(5294) when (flag_long='1') else '0';
	dataBufferOut(1571) <= dataBufferIn(6037) when (flag_long='1') else '0';
	dataBufferOut(1572) <= dataBufferIn( 636) when (flag_long='1') else '0';
	dataBufferOut(1573) <= dataBufferIn(1379) when (flag_long='1') else '0';
	dataBufferOut(1574) <= dataBufferIn(2122) when (flag_long='1') else '0';
	dataBufferOut(1575) <= dataBufferIn(2865) when (flag_long='1') else '0';
	dataBufferOut(1576) <= dataBufferIn(3608) when (flag_long='1') else '0';
	dataBufferOut(1577) <= dataBufferIn(4351) when (flag_long='1') else '0';
	dataBufferOut(1578) <= dataBufferIn(5094) when (flag_long='1') else '0';
	dataBufferOut(1579) <= dataBufferIn(5837) when (flag_long='1') else '0';
	dataBufferOut(1580) <= dataBufferIn( 436) when (flag_long='1') else '0';
	dataBufferOut(1581) <= dataBufferIn(1179) when (flag_long='1') else '0';
	dataBufferOut(1582) <= dataBufferIn(1922) when (flag_long='1') else '0';
	dataBufferOut(1583) <= dataBufferIn(2665) when (flag_long='1') else '0';
	dataBufferOut(1584) <= dataBufferIn(3408) when (flag_long='1') else '0';
	dataBufferOut(1585) <= dataBufferIn(4151) when (flag_long='1') else '0';
	dataBufferOut(1586) <= dataBufferIn(4894) when (flag_long='1') else '0';
	dataBufferOut(1587) <= dataBufferIn(5637) when (flag_long='1') else '0';
	dataBufferOut(1588) <= dataBufferIn( 236) when (flag_long='1') else '0';
	dataBufferOut(1589) <= dataBufferIn( 979) when (flag_long='1') else '0';
	dataBufferOut(1590) <= dataBufferIn(1722) when (flag_long='1') else '0';
	dataBufferOut(1591) <= dataBufferIn(2465) when (flag_long='1') else '0';
	dataBufferOut(1592) <= dataBufferIn(3208) when (flag_long='1') else '0';
	dataBufferOut(1593) <= dataBufferIn(3951) when (flag_long='1') else '0';
	dataBufferOut(1594) <= dataBufferIn(4694) when (flag_long='1') else '0';
	dataBufferOut(1595) <= dataBufferIn(5437) when (flag_long='1') else '0';
	dataBufferOut(1596) <= dataBufferIn(  36) when (flag_long='1') else '0';
	dataBufferOut(1597) <= dataBufferIn( 779) when (flag_long='1') else '0';
	dataBufferOut(1598) <= dataBufferIn(1522) when (flag_long='1') else '0';
	dataBufferOut(1599) <= dataBufferIn(2265) when (flag_long='1') else '0';
	dataBufferOut(1600) <= dataBufferIn(3008) when (flag_long='1') else '0';
	dataBufferOut(1601) <= dataBufferIn(3751) when (flag_long='1') else '0';
	dataBufferOut(1602) <= dataBufferIn(4494) when (flag_long='1') else '0';
	dataBufferOut(1603) <= dataBufferIn(5237) when (flag_long='1') else '0';
	dataBufferOut(1604) <= dataBufferIn(5980) when (flag_long='1') else '0';
	dataBufferOut(1605) <= dataBufferIn( 579) when (flag_long='1') else '0';
	dataBufferOut(1606) <= dataBufferIn(1322) when (flag_long='1') else '0';
	dataBufferOut(1607) <= dataBufferIn(2065) when (flag_long='1') else '0';
	dataBufferOut(1608) <= dataBufferIn(2808) when (flag_long='1') else '0';
	dataBufferOut(1609) <= dataBufferIn(3551) when (flag_long='1') else '0';
	dataBufferOut(1610) <= dataBufferIn(4294) when (flag_long='1') else '0';
	dataBufferOut(1611) <= dataBufferIn(5037) when (flag_long='1') else '0';
	dataBufferOut(1612) <= dataBufferIn(5780) when (flag_long='1') else '0';
	dataBufferOut(1613) <= dataBufferIn( 379) when (flag_long='1') else '0';
	dataBufferOut(1614) <= dataBufferIn(1122) when (flag_long='1') else '0';
	dataBufferOut(1615) <= dataBufferIn(1865) when (flag_long='1') else '0';
	dataBufferOut(1616) <= dataBufferIn(2608) when (flag_long='1') else '0';
	dataBufferOut(1617) <= dataBufferIn(3351) when (flag_long='1') else '0';
	dataBufferOut(1618) <= dataBufferIn(4094) when (flag_long='1') else '0';
	dataBufferOut(1619) <= dataBufferIn(4837) when (flag_long='1') else '0';
	dataBufferOut(1620) <= dataBufferIn(5580) when (flag_long='1') else '0';
	dataBufferOut(1621) <= dataBufferIn( 179) when (flag_long='1') else '0';
	dataBufferOut(1622) <= dataBufferIn( 922) when (flag_long='1') else '0';
	dataBufferOut(1623) <= dataBufferIn(1665) when (flag_long='1') else '0';
	dataBufferOut(1624) <= dataBufferIn(2408) when (flag_long='1') else '0';
	dataBufferOut(1625) <= dataBufferIn(3151) when (flag_long='1') else '0';
	dataBufferOut(1626) <= dataBufferIn(3894) when (flag_long='1') else '0';
	dataBufferOut(1627) <= dataBufferIn(4637) when (flag_long='1') else '0';
	dataBufferOut(1628) <= dataBufferIn(5380) when (flag_long='1') else '0';
	dataBufferOut(1629) <= dataBufferIn(6123) when (flag_long='1') else '0';
	dataBufferOut(1630) <= dataBufferIn( 722) when (flag_long='1') else '0';
	dataBufferOut(1631) <= dataBufferIn(1465) when (flag_long='1') else '0';
	dataBufferOut(1632) <= dataBufferIn(2208) when (flag_long='1') else '0';
	dataBufferOut(1633) <= dataBufferIn(2951) when (flag_long='1') else '0';
	dataBufferOut(1634) <= dataBufferIn(3694) when (flag_long='1') else '0';
	dataBufferOut(1635) <= dataBufferIn(4437) when (flag_long='1') else '0';
	dataBufferOut(1636) <= dataBufferIn(5180) when (flag_long='1') else '0';
	dataBufferOut(1637) <= dataBufferIn(5923) when (flag_long='1') else '0';
	dataBufferOut(1638) <= dataBufferIn( 522) when (flag_long='1') else '0';
	dataBufferOut(1639) <= dataBufferIn(1265) when (flag_long='1') else '0';
	dataBufferOut(1640) <= dataBufferIn(2008) when (flag_long='1') else '0';
	dataBufferOut(1641) <= dataBufferIn(2751) when (flag_long='1') else '0';
	dataBufferOut(1642) <= dataBufferIn(3494) when (flag_long='1') else '0';
	dataBufferOut(1643) <= dataBufferIn(4237) when (flag_long='1') else '0';
	dataBufferOut(1644) <= dataBufferIn(4980) when (flag_long='1') else '0';
	dataBufferOut(1645) <= dataBufferIn(5723) when (flag_long='1') else '0';
	dataBufferOut(1646) <= dataBufferIn( 322) when (flag_long='1') else '0';
	dataBufferOut(1647) <= dataBufferIn(1065) when (flag_long='1') else '0';
	dataBufferOut(1648) <= dataBufferIn(1808) when (flag_long='1') else '0';
	dataBufferOut(1649) <= dataBufferIn(2551) when (flag_long='1') else '0';
	dataBufferOut(1650) <= dataBufferIn(3294) when (flag_long='1') else '0';
	dataBufferOut(1651) <= dataBufferIn(4037) when (flag_long='1') else '0';
	dataBufferOut(1652) <= dataBufferIn(4780) when (flag_long='1') else '0';
	dataBufferOut(1653) <= dataBufferIn(5523) when (flag_long='1') else '0';
	dataBufferOut(1654) <= dataBufferIn( 122) when (flag_long='1') else '0';
	dataBufferOut(1655) <= dataBufferIn( 865) when (flag_long='1') else '0';
	dataBufferOut(1656) <= dataBufferIn(1608) when (flag_long='1') else '0';
	dataBufferOut(1657) <= dataBufferIn(2351) when (flag_long='1') else '0';
	dataBufferOut(1658) <= dataBufferIn(3094) when (flag_long='1') else '0';
	dataBufferOut(1659) <= dataBufferIn(3837) when (flag_long='1') else '0';
	dataBufferOut(1660) <= dataBufferIn(4580) when (flag_long='1') else '0';
	dataBufferOut(1661) <= dataBufferIn(5323) when (flag_long='1') else '0';
	dataBufferOut(1662) <= dataBufferIn(6066) when (flag_long='1') else '0';
	dataBufferOut(1663) <= dataBufferIn( 665) when (flag_long='1') else '0';
	dataBufferOut(1664) <= dataBufferIn(1408) when (flag_long='1') else '0';
	dataBufferOut(1665) <= dataBufferIn(2151) when (flag_long='1') else '0';
	dataBufferOut(1666) <= dataBufferIn(2894) when (flag_long='1') else '0';
	dataBufferOut(1667) <= dataBufferIn(3637) when (flag_long='1') else '0';
	dataBufferOut(1668) <= dataBufferIn(4380) when (flag_long='1') else '0';
	dataBufferOut(1669) <= dataBufferIn(5123) when (flag_long='1') else '0';
	dataBufferOut(1670) <= dataBufferIn(5866) when (flag_long='1') else '0';
	dataBufferOut(1671) <= dataBufferIn( 465) when (flag_long='1') else '0';
	dataBufferOut(1672) <= dataBufferIn(1208) when (flag_long='1') else '0';
	dataBufferOut(1673) <= dataBufferIn(1951) when (flag_long='1') else '0';
	dataBufferOut(1674) <= dataBufferIn(2694) when (flag_long='1') else '0';
	dataBufferOut(1675) <= dataBufferIn(3437) when (flag_long='1') else '0';
	dataBufferOut(1676) <= dataBufferIn(4180) when (flag_long='1') else '0';
	dataBufferOut(1677) <= dataBufferIn(4923) when (flag_long='1') else '0';
	dataBufferOut(1678) <= dataBufferIn(5666) when (flag_long='1') else '0';
	dataBufferOut(1679) <= dataBufferIn( 265) when (flag_long='1') else '0';
	dataBufferOut(1680) <= dataBufferIn(1008) when (flag_long='1') else '0';
	dataBufferOut(1681) <= dataBufferIn(1751) when (flag_long='1') else '0';
	dataBufferOut(1682) <= dataBufferIn(2494) when (flag_long='1') else '0';
	dataBufferOut(1683) <= dataBufferIn(3237) when (flag_long='1') else '0';
	dataBufferOut(1684) <= dataBufferIn(3980) when (flag_long='1') else '0';
	dataBufferOut(1685) <= dataBufferIn(4723) when (flag_long='1') else '0';
	dataBufferOut(1686) <= dataBufferIn(5466) when (flag_long='1') else '0';
	dataBufferOut(1687) <= dataBufferIn(  65) when (flag_long='1') else '0';
	dataBufferOut(1688) <= dataBufferIn( 808) when (flag_long='1') else '0';
	dataBufferOut(1689) <= dataBufferIn(1551) when (flag_long='1') else '0';
	dataBufferOut(1690) <= dataBufferIn(2294) when (flag_long='1') else '0';
	dataBufferOut(1691) <= dataBufferIn(3037) when (flag_long='1') else '0';
	dataBufferOut(1692) <= dataBufferIn(3780) when (flag_long='1') else '0';
	dataBufferOut(1693) <= dataBufferIn(4523) when (flag_long='1') else '0';
	dataBufferOut(1694) <= dataBufferIn(5266) when (flag_long='1') else '0';
	dataBufferOut(1695) <= dataBufferIn(6009) when (flag_long='1') else '0';
	dataBufferOut(1696) <= dataBufferIn( 608) when (flag_long='1') else '0';
	dataBufferOut(1697) <= dataBufferIn(1351) when (flag_long='1') else '0';
	dataBufferOut(1698) <= dataBufferIn(2094) when (flag_long='1') else '0';
	dataBufferOut(1699) <= dataBufferIn(2837) when (flag_long='1') else '0';
	dataBufferOut(1700) <= dataBufferIn(3580) when (flag_long='1') else '0';
	dataBufferOut(1701) <= dataBufferIn(4323) when (flag_long='1') else '0';
	dataBufferOut(1702) <= dataBufferIn(5066) when (flag_long='1') else '0';
	dataBufferOut(1703) <= dataBufferIn(5809) when (flag_long='1') else '0';
	dataBufferOut(1704) <= dataBufferIn( 408) when (flag_long='1') else '0';
	dataBufferOut(1705) <= dataBufferIn(1151) when (flag_long='1') else '0';
	dataBufferOut(1706) <= dataBufferIn(1894) when (flag_long='1') else '0';
	dataBufferOut(1707) <= dataBufferIn(2637) when (flag_long='1') else '0';
	dataBufferOut(1708) <= dataBufferIn(3380) when (flag_long='1') else '0';
	dataBufferOut(1709) <= dataBufferIn(4123) when (flag_long='1') else '0';
	dataBufferOut(1710) <= dataBufferIn(4866) when (flag_long='1') else '0';
	dataBufferOut(1711) <= dataBufferIn(5609) when (flag_long='1') else '0';
	dataBufferOut(1712) <= dataBufferIn( 208) when (flag_long='1') else '0';
	dataBufferOut(1713) <= dataBufferIn( 951) when (flag_long='1') else '0';
	dataBufferOut(1714) <= dataBufferIn(1694) when (flag_long='1') else '0';
	dataBufferOut(1715) <= dataBufferIn(2437) when (flag_long='1') else '0';
	dataBufferOut(1716) <= dataBufferIn(3180) when (flag_long='1') else '0';
	dataBufferOut(1717) <= dataBufferIn(3923) when (flag_long='1') else '0';
	dataBufferOut(1718) <= dataBufferIn(4666) when (flag_long='1') else '0';
	dataBufferOut(1719) <= dataBufferIn(5409) when (flag_long='1') else '0';
	dataBufferOut(1720) <= dataBufferIn(   8) when (flag_long='1') else '0';
	dataBufferOut(1721) <= dataBufferIn( 751) when (flag_long='1') else '0';
	dataBufferOut(1722) <= dataBufferIn(1494) when (flag_long='1') else '0';
	dataBufferOut(1723) <= dataBufferIn(2237) when (flag_long='1') else '0';
	dataBufferOut(1724) <= dataBufferIn(2980) when (flag_long='1') else '0';
	dataBufferOut(1725) <= dataBufferIn(3723) when (flag_long='1') else '0';
	dataBufferOut(1726) <= dataBufferIn(4466) when (flag_long='1') else '0';
	dataBufferOut(1727) <= dataBufferIn(5209) when (flag_long='1') else '0';
	dataBufferOut(1728) <= dataBufferIn(5952) when (flag_long='1') else '0';
	dataBufferOut(1729) <= dataBufferIn( 551) when (flag_long='1') else '0';
	dataBufferOut(1730) <= dataBufferIn(1294) when (flag_long='1') else '0';
	dataBufferOut(1731) <= dataBufferIn(2037) when (flag_long='1') else '0';
	dataBufferOut(1732) <= dataBufferIn(2780) when (flag_long='1') else '0';
	dataBufferOut(1733) <= dataBufferIn(3523) when (flag_long='1') else '0';
	dataBufferOut(1734) <= dataBufferIn(4266) when (flag_long='1') else '0';
	dataBufferOut(1735) <= dataBufferIn(5009) when (flag_long='1') else '0';
	dataBufferOut(1736) <= dataBufferIn(5752) when (flag_long='1') else '0';
	dataBufferOut(1737) <= dataBufferIn( 351) when (flag_long='1') else '0';
	dataBufferOut(1738) <= dataBufferIn(1094) when (flag_long='1') else '0';
	dataBufferOut(1739) <= dataBufferIn(1837) when (flag_long='1') else '0';
	dataBufferOut(1740) <= dataBufferIn(2580) when (flag_long='1') else '0';
	dataBufferOut(1741) <= dataBufferIn(3323) when (flag_long='1') else '0';
	dataBufferOut(1742) <= dataBufferIn(4066) when (flag_long='1') else '0';
	dataBufferOut(1743) <= dataBufferIn(4809) when (flag_long='1') else '0';
	dataBufferOut(1744) <= dataBufferIn(5552) when (flag_long='1') else '0';
	dataBufferOut(1745) <= dataBufferIn( 151) when (flag_long='1') else '0';
	dataBufferOut(1746) <= dataBufferIn( 894) when (flag_long='1') else '0';
	dataBufferOut(1747) <= dataBufferIn(1637) when (flag_long='1') else '0';
	dataBufferOut(1748) <= dataBufferIn(2380) when (flag_long='1') else '0';
	dataBufferOut(1749) <= dataBufferIn(3123) when (flag_long='1') else '0';
	dataBufferOut(1750) <= dataBufferIn(3866) when (flag_long='1') else '0';
	dataBufferOut(1751) <= dataBufferIn(4609) when (flag_long='1') else '0';
	dataBufferOut(1752) <= dataBufferIn(5352) when (flag_long='1') else '0';
	dataBufferOut(1753) <= dataBufferIn(6095) when (flag_long='1') else '0';
	dataBufferOut(1754) <= dataBufferIn( 694) when (flag_long='1') else '0';
	dataBufferOut(1755) <= dataBufferIn(1437) when (flag_long='1') else '0';
	dataBufferOut(1756) <= dataBufferIn(2180) when (flag_long='1') else '0';
	dataBufferOut(1757) <= dataBufferIn(2923) when (flag_long='1') else '0';
	dataBufferOut(1758) <= dataBufferIn(3666) when (flag_long='1') else '0';
	dataBufferOut(1759) <= dataBufferIn(4409) when (flag_long='1') else '0';
	dataBufferOut(1760) <= dataBufferIn(5152) when (flag_long='1') else '0';
	dataBufferOut(1761) <= dataBufferIn(5895) when (flag_long='1') else '0';
	dataBufferOut(1762) <= dataBufferIn( 494) when (flag_long='1') else '0';
	dataBufferOut(1763) <= dataBufferIn(1237) when (flag_long='1') else '0';
	dataBufferOut(1764) <= dataBufferIn(1980) when (flag_long='1') else '0';
	dataBufferOut(1765) <= dataBufferIn(2723) when (flag_long='1') else '0';
	dataBufferOut(1766) <= dataBufferIn(3466) when (flag_long='1') else '0';
	dataBufferOut(1767) <= dataBufferIn(4209) when (flag_long='1') else '0';
	dataBufferOut(1768) <= dataBufferIn(4952) when (flag_long='1') else '0';
	dataBufferOut(1769) <= dataBufferIn(5695) when (flag_long='1') else '0';
	dataBufferOut(1770) <= dataBufferIn( 294) when (flag_long='1') else '0';
	dataBufferOut(1771) <= dataBufferIn(1037) when (flag_long='1') else '0';
	dataBufferOut(1772) <= dataBufferIn(1780) when (flag_long='1') else '0';
	dataBufferOut(1773) <= dataBufferIn(2523) when (flag_long='1') else '0';
	dataBufferOut(1774) <= dataBufferIn(3266) when (flag_long='1') else '0';
	dataBufferOut(1775) <= dataBufferIn(4009) when (flag_long='1') else '0';
	dataBufferOut(1776) <= dataBufferIn(4752) when (flag_long='1') else '0';
	dataBufferOut(1777) <= dataBufferIn(5495) when (flag_long='1') else '0';
	dataBufferOut(1778) <= dataBufferIn(  94) when (flag_long='1') else '0';
	dataBufferOut(1779) <= dataBufferIn( 837) when (flag_long='1') else '0';
	dataBufferOut(1780) <= dataBufferIn(1580) when (flag_long='1') else '0';
	dataBufferOut(1781) <= dataBufferIn(2323) when (flag_long='1') else '0';
	dataBufferOut(1782) <= dataBufferIn(3066) when (flag_long='1') else '0';
	dataBufferOut(1783) <= dataBufferIn(3809) when (flag_long='1') else '0';
	dataBufferOut(1784) <= dataBufferIn(4552) when (flag_long='1') else '0';
	dataBufferOut(1785) <= dataBufferIn(5295) when (flag_long='1') else '0';
	dataBufferOut(1786) <= dataBufferIn(6038) when (flag_long='1') else '0';
	dataBufferOut(1787) <= dataBufferIn( 637) when (flag_long='1') else '0';
	dataBufferOut(1788) <= dataBufferIn(1380) when (flag_long='1') else '0';
	dataBufferOut(1789) <= dataBufferIn(2123) when (flag_long='1') else '0';
	dataBufferOut(1790) <= dataBufferIn(2866) when (flag_long='1') else '0';
	dataBufferOut(1791) <= dataBufferIn(3609) when (flag_long='1') else '0';
	dataBufferOut(1792) <= dataBufferIn(4352) when (flag_long='1') else '0';
	dataBufferOut(1793) <= dataBufferIn(5095) when (flag_long='1') else '0';
	dataBufferOut(1794) <= dataBufferIn(5838) when (flag_long='1') else '0';
	dataBufferOut(1795) <= dataBufferIn( 437) when (flag_long='1') else '0';
	dataBufferOut(1796) <= dataBufferIn(1180) when (flag_long='1') else '0';
	dataBufferOut(1797) <= dataBufferIn(1923) when (flag_long='1') else '0';
	dataBufferOut(1798) <= dataBufferIn(2666) when (flag_long='1') else '0';
	dataBufferOut(1799) <= dataBufferIn(3409) when (flag_long='1') else '0';
	dataBufferOut(1800) <= dataBufferIn(4152) when (flag_long='1') else '0';
	dataBufferOut(1801) <= dataBufferIn(4895) when (flag_long='1') else '0';
	dataBufferOut(1802) <= dataBufferIn(5638) when (flag_long='1') else '0';
	dataBufferOut(1803) <= dataBufferIn( 237) when (flag_long='1') else '0';
	dataBufferOut(1804) <= dataBufferIn( 980) when (flag_long='1') else '0';
	dataBufferOut(1805) <= dataBufferIn(1723) when (flag_long='1') else '0';
	dataBufferOut(1806) <= dataBufferIn(2466) when (flag_long='1') else '0';
	dataBufferOut(1807) <= dataBufferIn(3209) when (flag_long='1') else '0';
	dataBufferOut(1808) <= dataBufferIn(3952) when (flag_long='1') else '0';
	dataBufferOut(1809) <= dataBufferIn(4695) when (flag_long='1') else '0';
	dataBufferOut(1810) <= dataBufferIn(5438) when (flag_long='1') else '0';
	dataBufferOut(1811) <= dataBufferIn(  37) when (flag_long='1') else '0';
	dataBufferOut(1812) <= dataBufferIn( 780) when (flag_long='1') else '0';
	dataBufferOut(1813) <= dataBufferIn(1523) when (flag_long='1') else '0';
	dataBufferOut(1814) <= dataBufferIn(2266) when (flag_long='1') else '0';
	dataBufferOut(1815) <= dataBufferIn(3009) when (flag_long='1') else '0';
	dataBufferOut(1816) <= dataBufferIn(3752) when (flag_long='1') else '0';
	dataBufferOut(1817) <= dataBufferIn(4495) when (flag_long='1') else '0';
	dataBufferOut(1818) <= dataBufferIn(5238) when (flag_long='1') else '0';
	dataBufferOut(1819) <= dataBufferIn(5981) when (flag_long='1') else '0';
	dataBufferOut(1820) <= dataBufferIn( 580) when (flag_long='1') else '0';
	dataBufferOut(1821) <= dataBufferIn(1323) when (flag_long='1') else '0';
	dataBufferOut(1822) <= dataBufferIn(2066) when (flag_long='1') else '0';
	dataBufferOut(1823) <= dataBufferIn(2809) when (flag_long='1') else '0';
	dataBufferOut(1824) <= dataBufferIn(3552) when (flag_long='1') else '0';
	dataBufferOut(1825) <= dataBufferIn(4295) when (flag_long='1') else '0';
	dataBufferOut(1826) <= dataBufferIn(5038) when (flag_long='1') else '0';
	dataBufferOut(1827) <= dataBufferIn(5781) when (flag_long='1') else '0';
	dataBufferOut(1828) <= dataBufferIn( 380) when (flag_long='1') else '0';
	dataBufferOut(1829) <= dataBufferIn(1123) when (flag_long='1') else '0';
	dataBufferOut(1830) <= dataBufferIn(1866) when (flag_long='1') else '0';
	dataBufferOut(1831) <= dataBufferIn(2609) when (flag_long='1') else '0';
	dataBufferOut(1832) <= dataBufferIn(3352) when (flag_long='1') else '0';
	dataBufferOut(1833) <= dataBufferIn(4095) when (flag_long='1') else '0';
	dataBufferOut(1834) <= dataBufferIn(4838) when (flag_long='1') else '0';
	dataBufferOut(1835) <= dataBufferIn(5581) when (flag_long='1') else '0';
	dataBufferOut(1836) <= dataBufferIn( 180) when (flag_long='1') else '0';
	dataBufferOut(1837) <= dataBufferIn( 923) when (flag_long='1') else '0';
	dataBufferOut(1838) <= dataBufferIn(1666) when (flag_long='1') else '0';
	dataBufferOut(1839) <= dataBufferIn(2409) when (flag_long='1') else '0';
	dataBufferOut(1840) <= dataBufferIn(3152) when (flag_long='1') else '0';
	dataBufferOut(1841) <= dataBufferIn(3895) when (flag_long='1') else '0';
	dataBufferOut(1842) <= dataBufferIn(4638) when (flag_long='1') else '0';
	dataBufferOut(1843) <= dataBufferIn(5381) when (flag_long='1') else '0';
	dataBufferOut(1844) <= dataBufferIn(6124) when (flag_long='1') else '0';
	dataBufferOut(1845) <= dataBufferIn( 723) when (flag_long='1') else '0';
	dataBufferOut(1846) <= dataBufferIn(1466) when (flag_long='1') else '0';
	dataBufferOut(1847) <= dataBufferIn(2209) when (flag_long='1') else '0';
	dataBufferOut(1848) <= dataBufferIn(2952) when (flag_long='1') else '0';
	dataBufferOut(1849) <= dataBufferIn(3695) when (flag_long='1') else '0';
	dataBufferOut(1850) <= dataBufferIn(4438) when (flag_long='1') else '0';
	dataBufferOut(1851) <= dataBufferIn(5181) when (flag_long='1') else '0';
	dataBufferOut(1852) <= dataBufferIn(5924) when (flag_long='1') else '0';
	dataBufferOut(1853) <= dataBufferIn( 523) when (flag_long='1') else '0';
	dataBufferOut(1854) <= dataBufferIn(1266) when (flag_long='1') else '0';
	dataBufferOut(1855) <= dataBufferIn(2009) when (flag_long='1') else '0';
	dataBufferOut(1856) <= dataBufferIn(2752) when (flag_long='1') else '0';
	dataBufferOut(1857) <= dataBufferIn(3495) when (flag_long='1') else '0';
	dataBufferOut(1858) <= dataBufferIn(4238) when (flag_long='1') else '0';
	dataBufferOut(1859) <= dataBufferIn(4981) when (flag_long='1') else '0';
	dataBufferOut(1860) <= dataBufferIn(5724) when (flag_long='1') else '0';
	dataBufferOut(1861) <= dataBufferIn( 323) when (flag_long='1') else '0';
	dataBufferOut(1862) <= dataBufferIn(1066) when (flag_long='1') else '0';
	dataBufferOut(1863) <= dataBufferIn(1809) when (flag_long='1') else '0';
	dataBufferOut(1864) <= dataBufferIn(2552) when (flag_long='1') else '0';
	dataBufferOut(1865) <= dataBufferIn(3295) when (flag_long='1') else '0';
	dataBufferOut(1866) <= dataBufferIn(4038) when (flag_long='1') else '0';
	dataBufferOut(1867) <= dataBufferIn(4781) when (flag_long='1') else '0';
	dataBufferOut(1868) <= dataBufferIn(5524) when (flag_long='1') else '0';
	dataBufferOut(1869) <= dataBufferIn( 123) when (flag_long='1') else '0';
	dataBufferOut(1870) <= dataBufferIn( 866) when (flag_long='1') else '0';
	dataBufferOut(1871) <= dataBufferIn(1609) when (flag_long='1') else '0';
	dataBufferOut(1872) <= dataBufferIn(2352) when (flag_long='1') else '0';
	dataBufferOut(1873) <= dataBufferIn(3095) when (flag_long='1') else '0';
	dataBufferOut(1874) <= dataBufferIn(3838) when (flag_long='1') else '0';
	dataBufferOut(1875) <= dataBufferIn(4581) when (flag_long='1') else '0';
	dataBufferOut(1876) <= dataBufferIn(5324) when (flag_long='1') else '0';
	dataBufferOut(1877) <= dataBufferIn(6067) when (flag_long='1') else '0';
	dataBufferOut(1878) <= dataBufferIn( 666) when (flag_long='1') else '0';
	dataBufferOut(1879) <= dataBufferIn(1409) when (flag_long='1') else '0';
	dataBufferOut(1880) <= dataBufferIn(2152) when (flag_long='1') else '0';
	dataBufferOut(1881) <= dataBufferIn(2895) when (flag_long='1') else '0';
	dataBufferOut(1882) <= dataBufferIn(3638) when (flag_long='1') else '0';
	dataBufferOut(1883) <= dataBufferIn(4381) when (flag_long='1') else '0';
	dataBufferOut(1884) <= dataBufferIn(5124) when (flag_long='1') else '0';
	dataBufferOut(1885) <= dataBufferIn(5867) when (flag_long='1') else '0';
	dataBufferOut(1886) <= dataBufferIn( 466) when (flag_long='1') else '0';
	dataBufferOut(1887) <= dataBufferIn(1209) when (flag_long='1') else '0';
	dataBufferOut(1888) <= dataBufferIn(1952) when (flag_long='1') else '0';
	dataBufferOut(1889) <= dataBufferIn(2695) when (flag_long='1') else '0';
	dataBufferOut(1890) <= dataBufferIn(3438) when (flag_long='1') else '0';
	dataBufferOut(1891) <= dataBufferIn(4181) when (flag_long='1') else '0';
	dataBufferOut(1892) <= dataBufferIn(4924) when (flag_long='1') else '0';
	dataBufferOut(1893) <= dataBufferIn(5667) when (flag_long='1') else '0';
	dataBufferOut(1894) <= dataBufferIn( 266) when (flag_long='1') else '0';
	dataBufferOut(1895) <= dataBufferIn(1009) when (flag_long='1') else '0';
	dataBufferOut(1896) <= dataBufferIn(1752) when (flag_long='1') else '0';
	dataBufferOut(1897) <= dataBufferIn(2495) when (flag_long='1') else '0';
	dataBufferOut(1898) <= dataBufferIn(3238) when (flag_long='1') else '0';
	dataBufferOut(1899) <= dataBufferIn(3981) when (flag_long='1') else '0';
	dataBufferOut(1900) <= dataBufferIn(4724) when (flag_long='1') else '0';
	dataBufferOut(1901) <= dataBufferIn(5467) when (flag_long='1') else '0';
	dataBufferOut(1902) <= dataBufferIn(  66) when (flag_long='1') else '0';
	dataBufferOut(1903) <= dataBufferIn( 809) when (flag_long='1') else '0';
	dataBufferOut(1904) <= dataBufferIn(1552) when (flag_long='1') else '0';
	dataBufferOut(1905) <= dataBufferIn(2295) when (flag_long='1') else '0';
	dataBufferOut(1906) <= dataBufferIn(3038) when (flag_long='1') else '0';
	dataBufferOut(1907) <= dataBufferIn(3781) when (flag_long='1') else '0';
	dataBufferOut(1908) <= dataBufferIn(4524) when (flag_long='1') else '0';
	dataBufferOut(1909) <= dataBufferIn(5267) when (flag_long='1') else '0';
	dataBufferOut(1910) <= dataBufferIn(6010) when (flag_long='1') else '0';
	dataBufferOut(1911) <= dataBufferIn( 609) when (flag_long='1') else '0';
	dataBufferOut(1912) <= dataBufferIn(1352) when (flag_long='1') else '0';
	dataBufferOut(1913) <= dataBufferIn(2095) when (flag_long='1') else '0';
	dataBufferOut(1914) <= dataBufferIn(2838) when (flag_long='1') else '0';
	dataBufferOut(1915) <= dataBufferIn(3581) when (flag_long='1') else '0';
	dataBufferOut(1916) <= dataBufferIn(4324) when (flag_long='1') else '0';
	dataBufferOut(1917) <= dataBufferIn(5067) when (flag_long='1') else '0';
	dataBufferOut(1918) <= dataBufferIn(5810) when (flag_long='1') else '0';
	dataBufferOut(1919) <= dataBufferIn( 409) when (flag_long='1') else '0';
	dataBufferOut(1920) <= dataBufferIn(1152) when (flag_long='1') else '0';
	dataBufferOut(1921) <= dataBufferIn(1895) when (flag_long='1') else '0';
	dataBufferOut(1922) <= dataBufferIn(2638) when (flag_long='1') else '0';
	dataBufferOut(1923) <= dataBufferIn(3381) when (flag_long='1') else '0';
	dataBufferOut(1924) <= dataBufferIn(4124) when (flag_long='1') else '0';
	dataBufferOut(1925) <= dataBufferIn(4867) when (flag_long='1') else '0';
	dataBufferOut(1926) <= dataBufferIn(5610) when (flag_long='1') else '0';
	dataBufferOut(1927) <= dataBufferIn( 209) when (flag_long='1') else '0';
	dataBufferOut(1928) <= dataBufferIn( 952) when (flag_long='1') else '0';
	dataBufferOut(1929) <= dataBufferIn(1695) when (flag_long='1') else '0';
	dataBufferOut(1930) <= dataBufferIn(2438) when (flag_long='1') else '0';
	dataBufferOut(1931) <= dataBufferIn(3181) when (flag_long='1') else '0';
	dataBufferOut(1932) <= dataBufferIn(3924) when (flag_long='1') else '0';
	dataBufferOut(1933) <= dataBufferIn(4667) when (flag_long='1') else '0';
	dataBufferOut(1934) <= dataBufferIn(5410) when (flag_long='1') else '0';
	dataBufferOut(1935) <= dataBufferIn(   9) when (flag_long='1') else '0';
	dataBufferOut(1936) <= dataBufferIn( 752) when (flag_long='1') else '0';
	dataBufferOut(1937) <= dataBufferIn(1495) when (flag_long='1') else '0';
	dataBufferOut(1938) <= dataBufferIn(2238) when (flag_long='1') else '0';
	dataBufferOut(1939) <= dataBufferIn(2981) when (flag_long='1') else '0';
	dataBufferOut(1940) <= dataBufferIn(3724) when (flag_long='1') else '0';
	dataBufferOut(1941) <= dataBufferIn(4467) when (flag_long='1') else '0';
	dataBufferOut(1942) <= dataBufferIn(5210) when (flag_long='1') else '0';
	dataBufferOut(1943) <= dataBufferIn(5953) when (flag_long='1') else '0';
	dataBufferOut(1944) <= dataBufferIn( 552) when (flag_long='1') else '0';
	dataBufferOut(1945) <= dataBufferIn(1295) when (flag_long='1') else '0';
	dataBufferOut(1946) <= dataBufferIn(2038) when (flag_long='1') else '0';
	dataBufferOut(1947) <= dataBufferIn(2781) when (flag_long='1') else '0';
	dataBufferOut(1948) <= dataBufferIn(3524) when (flag_long='1') else '0';
	dataBufferOut(1949) <= dataBufferIn(4267) when (flag_long='1') else '0';
	dataBufferOut(1950) <= dataBufferIn(5010) when (flag_long='1') else '0';
	dataBufferOut(1951) <= dataBufferIn(5753) when (flag_long='1') else '0';
	dataBufferOut(1952) <= dataBufferIn( 352) when (flag_long='1') else '0';
	dataBufferOut(1953) <= dataBufferIn(1095) when (flag_long='1') else '0';
	dataBufferOut(1954) <= dataBufferIn(1838) when (flag_long='1') else '0';
	dataBufferOut(1955) <= dataBufferIn(2581) when (flag_long='1') else '0';
	dataBufferOut(1956) <= dataBufferIn(3324) when (flag_long='1') else '0';
	dataBufferOut(1957) <= dataBufferIn(4067) when (flag_long='1') else '0';
	dataBufferOut(1958) <= dataBufferIn(4810) when (flag_long='1') else '0';
	dataBufferOut(1959) <= dataBufferIn(5553) when (flag_long='1') else '0';
	dataBufferOut(1960) <= dataBufferIn( 152) when (flag_long='1') else '0';
	dataBufferOut(1961) <= dataBufferIn( 895) when (flag_long='1') else '0';
	dataBufferOut(1962) <= dataBufferIn(1638) when (flag_long='1') else '0';
	dataBufferOut(1963) <= dataBufferIn(2381) when (flag_long='1') else '0';
	dataBufferOut(1964) <= dataBufferIn(3124) when (flag_long='1') else '0';
	dataBufferOut(1965) <= dataBufferIn(3867) when (flag_long='1') else '0';
	dataBufferOut(1966) <= dataBufferIn(4610) when (flag_long='1') else '0';
	dataBufferOut(1967) <= dataBufferIn(5353) when (flag_long='1') else '0';
	dataBufferOut(1968) <= dataBufferIn(6096) when (flag_long='1') else '0';
	dataBufferOut(1969) <= dataBufferIn( 695) when (flag_long='1') else '0';
	dataBufferOut(1970) <= dataBufferIn(1438) when (flag_long='1') else '0';
	dataBufferOut(1971) <= dataBufferIn(2181) when (flag_long='1') else '0';
	dataBufferOut(1972) <= dataBufferIn(2924) when (flag_long='1') else '0';
	dataBufferOut(1973) <= dataBufferIn(3667) when (flag_long='1') else '0';
	dataBufferOut(1974) <= dataBufferIn(4410) when (flag_long='1') else '0';
	dataBufferOut(1975) <= dataBufferIn(5153) when (flag_long='1') else '0';
	dataBufferOut(1976) <= dataBufferIn(5896) when (flag_long='1') else '0';
	dataBufferOut(1977) <= dataBufferIn( 495) when (flag_long='1') else '0';
	dataBufferOut(1978) <= dataBufferIn(1238) when (flag_long='1') else '0';
	dataBufferOut(1979) <= dataBufferIn(1981) when (flag_long='1') else '0';
	dataBufferOut(1980) <= dataBufferIn(2724) when (flag_long='1') else '0';
	dataBufferOut(1981) <= dataBufferIn(3467) when (flag_long='1') else '0';
	dataBufferOut(1982) <= dataBufferIn(4210) when (flag_long='1') else '0';
	dataBufferOut(1983) <= dataBufferIn(4953) when (flag_long='1') else '0';
	dataBufferOut(1984) <= dataBufferIn(5696) when (flag_long='1') else '0';
	dataBufferOut(1985) <= dataBufferIn( 295) when (flag_long='1') else '0';
	dataBufferOut(1986) <= dataBufferIn(1038) when (flag_long='1') else '0';
	dataBufferOut(1987) <= dataBufferIn(1781) when (flag_long='1') else '0';
	dataBufferOut(1988) <= dataBufferIn(2524) when (flag_long='1') else '0';
	dataBufferOut(1989) <= dataBufferIn(3267) when (flag_long='1') else '0';
	dataBufferOut(1990) <= dataBufferIn(4010) when (flag_long='1') else '0';
	dataBufferOut(1991) <= dataBufferIn(4753) when (flag_long='1') else '0';
	dataBufferOut(1992) <= dataBufferIn(5496) when (flag_long='1') else '0';
	dataBufferOut(1993) <= dataBufferIn(  95) when (flag_long='1') else '0';
	dataBufferOut(1994) <= dataBufferIn( 838) when (flag_long='1') else '0';
	dataBufferOut(1995) <= dataBufferIn(1581) when (flag_long='1') else '0';
	dataBufferOut(1996) <= dataBufferIn(2324) when (flag_long='1') else '0';
	dataBufferOut(1997) <= dataBufferIn(3067) when (flag_long='1') else '0';
	dataBufferOut(1998) <= dataBufferIn(3810) when (flag_long='1') else '0';
	dataBufferOut(1999) <= dataBufferIn(4553) when (flag_long='1') else '0';
	dataBufferOut(2000) <= dataBufferIn(5296) when (flag_long='1') else '0';
	dataBufferOut(2001) <= dataBufferIn(6039) when (flag_long='1') else '0';
	dataBufferOut(2002) <= dataBufferIn( 638) when (flag_long='1') else '0';
	dataBufferOut(2003) <= dataBufferIn(1381) when (flag_long='1') else '0';
	dataBufferOut(2004) <= dataBufferIn(2124) when (flag_long='1') else '0';
	dataBufferOut(2005) <= dataBufferIn(2867) when (flag_long='1') else '0';
	dataBufferOut(2006) <= dataBufferIn(3610) when (flag_long='1') else '0';
	dataBufferOut(2007) <= dataBufferIn(4353) when (flag_long='1') else '0';
	dataBufferOut(2008) <= dataBufferIn(5096) when (flag_long='1') else '0';
	dataBufferOut(2009) <= dataBufferIn(5839) when (flag_long='1') else '0';
	dataBufferOut(2010) <= dataBufferIn( 438) when (flag_long='1') else '0';
	dataBufferOut(2011) <= dataBufferIn(1181) when (flag_long='1') else '0';
	dataBufferOut(2012) <= dataBufferIn(1924) when (flag_long='1') else '0';
	dataBufferOut(2013) <= dataBufferIn(2667) when (flag_long='1') else '0';
	dataBufferOut(2014) <= dataBufferIn(3410) when (flag_long='1') else '0';
	dataBufferOut(2015) <= dataBufferIn(4153) when (flag_long='1') else '0';
	dataBufferOut(2016) <= dataBufferIn(4896) when (flag_long='1') else '0';
	dataBufferOut(2017) <= dataBufferIn(5639) when (flag_long='1') else '0';
	dataBufferOut(2018) <= dataBufferIn( 238) when (flag_long='1') else '0';
	dataBufferOut(2019) <= dataBufferIn( 981) when (flag_long='1') else '0';
	dataBufferOut(2020) <= dataBufferIn(1724) when (flag_long='1') else '0';
	dataBufferOut(2021) <= dataBufferIn(2467) when (flag_long='1') else '0';
	dataBufferOut(2022) <= dataBufferIn(3210) when (flag_long='1') else '0';
	dataBufferOut(2023) <= dataBufferIn(3953) when (flag_long='1') else '0';
	dataBufferOut(2024) <= dataBufferIn(4696) when (flag_long='1') else '0';
	dataBufferOut(2025) <= dataBufferIn(5439) when (flag_long='1') else '0';
	dataBufferOut(2026) <= dataBufferIn(  38) when (flag_long='1') else '0';
	dataBufferOut(2027) <= dataBufferIn( 781) when (flag_long='1') else '0';
	dataBufferOut(2028) <= dataBufferIn(1524) when (flag_long='1') else '0';
	dataBufferOut(2029) <= dataBufferIn(2267) when (flag_long='1') else '0';
	dataBufferOut(2030) <= dataBufferIn(3010) when (flag_long='1') else '0';
	dataBufferOut(2031) <= dataBufferIn(3753) when (flag_long='1') else '0';
	dataBufferOut(2032) <= dataBufferIn(4496) when (flag_long='1') else '0';
	dataBufferOut(2033) <= dataBufferIn(5239) when (flag_long='1') else '0';
	dataBufferOut(2034) <= dataBufferIn(5982) when (flag_long='1') else '0';
	dataBufferOut(2035) <= dataBufferIn( 581) when (flag_long='1') else '0';
	dataBufferOut(2036) <= dataBufferIn(1324) when (flag_long='1') else '0';
	dataBufferOut(2037) <= dataBufferIn(2067) when (flag_long='1') else '0';
	dataBufferOut(2038) <= dataBufferIn(2810) when (flag_long='1') else '0';
	dataBufferOut(2039) <= dataBufferIn(3553) when (flag_long='1') else '0';
	dataBufferOut(2040) <= dataBufferIn(4296) when (flag_long='1') else '0';
	dataBufferOut(2041) <= dataBufferIn(5039) when (flag_long='1') else '0';
	dataBufferOut(2042) <= dataBufferIn(5782) when (flag_long='1') else '0';
	dataBufferOut(2043) <= dataBufferIn( 381) when (flag_long='1') else '0';
	dataBufferOut(2044) <= dataBufferIn(1124) when (flag_long='1') else '0';
	dataBufferOut(2045) <= dataBufferIn(1867) when (flag_long='1') else '0';
	dataBufferOut(2046) <= dataBufferIn(2610) when (flag_long='1') else '0';
	dataBufferOut(2047) <= dataBufferIn(3353) when (flag_long='1') else '0';
	dataBufferOut(2048) <= dataBufferIn(4096) when (flag_long='1') else '0';
	dataBufferOut(2049) <= dataBufferIn(4839) when (flag_long='1') else '0';
	dataBufferOut(2050) <= dataBufferIn(5582) when (flag_long='1') else '0';
	dataBufferOut(2051) <= dataBufferIn( 181) when (flag_long='1') else '0';
	dataBufferOut(2052) <= dataBufferIn( 924) when (flag_long='1') else '0';
	dataBufferOut(2053) <= dataBufferIn(1667) when (flag_long='1') else '0';
	dataBufferOut(2054) <= dataBufferIn(2410) when (flag_long='1') else '0';
	dataBufferOut(2055) <= dataBufferIn(3153) when (flag_long='1') else '0';
	dataBufferOut(2056) <= dataBufferIn(3896) when (flag_long='1') else '0';
	dataBufferOut(2057) <= dataBufferIn(4639) when (flag_long='1') else '0';
	dataBufferOut(2058) <= dataBufferIn(5382) when (flag_long='1') else '0';
	dataBufferOut(2059) <= dataBufferIn(6125) when (flag_long='1') else '0';
	dataBufferOut(2060) <= dataBufferIn( 724) when (flag_long='1') else '0';
	dataBufferOut(2061) <= dataBufferIn(1467) when (flag_long='1') else '0';
	dataBufferOut(2062) <= dataBufferIn(2210) when (flag_long='1') else '0';
	dataBufferOut(2063) <= dataBufferIn(2953) when (flag_long='1') else '0';
	dataBufferOut(2064) <= dataBufferIn(3696) when (flag_long='1') else '0';
	dataBufferOut(2065) <= dataBufferIn(4439) when (flag_long='1') else '0';
	dataBufferOut(2066) <= dataBufferIn(5182) when (flag_long='1') else '0';
	dataBufferOut(2067) <= dataBufferIn(5925) when (flag_long='1') else '0';
	dataBufferOut(2068) <= dataBufferIn( 524) when (flag_long='1') else '0';
	dataBufferOut(2069) <= dataBufferIn(1267) when (flag_long='1') else '0';
	dataBufferOut(2070) <= dataBufferIn(2010) when (flag_long='1') else '0';
	dataBufferOut(2071) <= dataBufferIn(2753) when (flag_long='1') else '0';
	dataBufferOut(2072) <= dataBufferIn(3496) when (flag_long='1') else '0';
	dataBufferOut(2073) <= dataBufferIn(4239) when (flag_long='1') else '0';
	dataBufferOut(2074) <= dataBufferIn(4982) when (flag_long='1') else '0';
	dataBufferOut(2075) <= dataBufferIn(5725) when (flag_long='1') else '0';
	dataBufferOut(2076) <= dataBufferIn( 324) when (flag_long='1') else '0';
	dataBufferOut(2077) <= dataBufferIn(1067) when (flag_long='1') else '0';
	dataBufferOut(2078) <= dataBufferIn(1810) when (flag_long='1') else '0';
	dataBufferOut(2079) <= dataBufferIn(2553) when (flag_long='1') else '0';
	dataBufferOut(2080) <= dataBufferIn(3296) when (flag_long='1') else '0';
	dataBufferOut(2081) <= dataBufferIn(4039) when (flag_long='1') else '0';
	dataBufferOut(2082) <= dataBufferIn(4782) when (flag_long='1') else '0';
	dataBufferOut(2083) <= dataBufferIn(5525) when (flag_long='1') else '0';
	dataBufferOut(2084) <= dataBufferIn( 124) when (flag_long='1') else '0';
	dataBufferOut(2085) <= dataBufferIn( 867) when (flag_long='1') else '0';
	dataBufferOut(2086) <= dataBufferIn(1610) when (flag_long='1') else '0';
	dataBufferOut(2087) <= dataBufferIn(2353) when (flag_long='1') else '0';
	dataBufferOut(2088) <= dataBufferIn(3096) when (flag_long='1') else '0';
	dataBufferOut(2089) <= dataBufferIn(3839) when (flag_long='1') else '0';
	dataBufferOut(2090) <= dataBufferIn(4582) when (flag_long='1') else '0';
	dataBufferOut(2091) <= dataBufferIn(5325) when (flag_long='1') else '0';
	dataBufferOut(2092) <= dataBufferIn(6068) when (flag_long='1') else '0';
	dataBufferOut(2093) <= dataBufferIn( 667) when (flag_long='1') else '0';
	dataBufferOut(2094) <= dataBufferIn(1410) when (flag_long='1') else '0';
	dataBufferOut(2095) <= dataBufferIn(2153) when (flag_long='1') else '0';
	dataBufferOut(2096) <= dataBufferIn(2896) when (flag_long='1') else '0';
	dataBufferOut(2097) <= dataBufferIn(3639) when (flag_long='1') else '0';
	dataBufferOut(2098) <= dataBufferIn(4382) when (flag_long='1') else '0';
	dataBufferOut(2099) <= dataBufferIn(5125) when (flag_long='1') else '0';
	dataBufferOut(2100) <= dataBufferIn(5868) when (flag_long='1') else '0';
	dataBufferOut(2101) <= dataBufferIn( 467) when (flag_long='1') else '0';
	dataBufferOut(2102) <= dataBufferIn(1210) when (flag_long='1') else '0';
	dataBufferOut(2103) <= dataBufferIn(1953) when (flag_long='1') else '0';
	dataBufferOut(2104) <= dataBufferIn(2696) when (flag_long='1') else '0';
	dataBufferOut(2105) <= dataBufferIn(3439) when (flag_long='1') else '0';
	dataBufferOut(2106) <= dataBufferIn(4182) when (flag_long='1') else '0';
	dataBufferOut(2107) <= dataBufferIn(4925) when (flag_long='1') else '0';
	dataBufferOut(2108) <= dataBufferIn(5668) when (flag_long='1') else '0';
	dataBufferOut(2109) <= dataBufferIn( 267) when (flag_long='1') else '0';
	dataBufferOut(2110) <= dataBufferIn(1010) when (flag_long='1') else '0';
	dataBufferOut(2111) <= dataBufferIn(1753) when (flag_long='1') else '0';
	dataBufferOut(2112) <= dataBufferIn(2496) when (flag_long='1') else '0';
	dataBufferOut(2113) <= dataBufferIn(3239) when (flag_long='1') else '0';
	dataBufferOut(2114) <= dataBufferIn(3982) when (flag_long='1') else '0';
	dataBufferOut(2115) <= dataBufferIn(4725) when (flag_long='1') else '0';
	dataBufferOut(2116) <= dataBufferIn(5468) when (flag_long='1') else '0';
	dataBufferOut(2117) <= dataBufferIn(  67) when (flag_long='1') else '0';
	dataBufferOut(2118) <= dataBufferIn( 810) when (flag_long='1') else '0';
	dataBufferOut(2119) <= dataBufferIn(1553) when (flag_long='1') else '0';
	dataBufferOut(2120) <= dataBufferIn(2296) when (flag_long='1') else '0';
	dataBufferOut(2121) <= dataBufferIn(3039) when (flag_long='1') else '0';
	dataBufferOut(2122) <= dataBufferIn(3782) when (flag_long='1') else '0';
	dataBufferOut(2123) <= dataBufferIn(4525) when (flag_long='1') else '0';
	dataBufferOut(2124) <= dataBufferIn(5268) when (flag_long='1') else '0';
	dataBufferOut(2125) <= dataBufferIn(6011) when (flag_long='1') else '0';
	dataBufferOut(2126) <= dataBufferIn( 610) when (flag_long='1') else '0';
	dataBufferOut(2127) <= dataBufferIn(1353) when (flag_long='1') else '0';
	dataBufferOut(2128) <= dataBufferIn(2096) when (flag_long='1') else '0';
	dataBufferOut(2129) <= dataBufferIn(2839) when (flag_long='1') else '0';
	dataBufferOut(2130) <= dataBufferIn(3582) when (flag_long='1') else '0';
	dataBufferOut(2131) <= dataBufferIn(4325) when (flag_long='1') else '0';
	dataBufferOut(2132) <= dataBufferIn(5068) when (flag_long='1') else '0';
	dataBufferOut(2133) <= dataBufferIn(5811) when (flag_long='1') else '0';
	dataBufferOut(2134) <= dataBufferIn( 410) when (flag_long='1') else '0';
	dataBufferOut(2135) <= dataBufferIn(1153) when (flag_long='1') else '0';
	dataBufferOut(2136) <= dataBufferIn(1896) when (flag_long='1') else '0';
	dataBufferOut(2137) <= dataBufferIn(2639) when (flag_long='1') else '0';
	dataBufferOut(2138) <= dataBufferIn(3382) when (flag_long='1') else '0';
	dataBufferOut(2139) <= dataBufferIn(4125) when (flag_long='1') else '0';
	dataBufferOut(2140) <= dataBufferIn(4868) when (flag_long='1') else '0';
	dataBufferOut(2141) <= dataBufferIn(5611) when (flag_long='1') else '0';
	dataBufferOut(2142) <= dataBufferIn( 210) when (flag_long='1') else '0';
	dataBufferOut(2143) <= dataBufferIn( 953) when (flag_long='1') else '0';
	dataBufferOut(2144) <= dataBufferIn(1696) when (flag_long='1') else '0';
	dataBufferOut(2145) <= dataBufferIn(2439) when (flag_long='1') else '0';
	dataBufferOut(2146) <= dataBufferIn(3182) when (flag_long='1') else '0';
	dataBufferOut(2147) <= dataBufferIn(3925) when (flag_long='1') else '0';
	dataBufferOut(2148) <= dataBufferIn(4668) when (flag_long='1') else '0';
	dataBufferOut(2149) <= dataBufferIn(5411) when (flag_long='1') else '0';
	dataBufferOut(2150) <= dataBufferIn(  10) when (flag_long='1') else '0';
	dataBufferOut(2151) <= dataBufferIn( 753) when (flag_long='1') else '0';
	dataBufferOut(2152) <= dataBufferIn(1496) when (flag_long='1') else '0';
	dataBufferOut(2153) <= dataBufferIn(2239) when (flag_long='1') else '0';
	dataBufferOut(2154) <= dataBufferIn(2982) when (flag_long='1') else '0';
	dataBufferOut(2155) <= dataBufferIn(3725) when (flag_long='1') else '0';
	dataBufferOut(2156) <= dataBufferIn(4468) when (flag_long='1') else '0';
	dataBufferOut(2157) <= dataBufferIn(5211) when (flag_long='1') else '0';
	dataBufferOut(2158) <= dataBufferIn(5954) when (flag_long='1') else '0';
	dataBufferOut(2159) <= dataBufferIn( 553) when (flag_long='1') else '0';
	dataBufferOut(2160) <= dataBufferIn(1296) when (flag_long='1') else '0';
	dataBufferOut(2161) <= dataBufferIn(2039) when (flag_long='1') else '0';
	dataBufferOut(2162) <= dataBufferIn(2782) when (flag_long='1') else '0';
	dataBufferOut(2163) <= dataBufferIn(3525) when (flag_long='1') else '0';
	dataBufferOut(2164) <= dataBufferIn(4268) when (flag_long='1') else '0';
	dataBufferOut(2165) <= dataBufferIn(5011) when (flag_long='1') else '0';
	dataBufferOut(2166) <= dataBufferIn(5754) when (flag_long='1') else '0';
	dataBufferOut(2167) <= dataBufferIn( 353) when (flag_long='1') else '0';
	dataBufferOut(2168) <= dataBufferIn(1096) when (flag_long='1') else '0';
	dataBufferOut(2169) <= dataBufferIn(1839) when (flag_long='1') else '0';
	dataBufferOut(2170) <= dataBufferIn(2582) when (flag_long='1') else '0';
	dataBufferOut(2171) <= dataBufferIn(3325) when (flag_long='1') else '0';
	dataBufferOut(2172) <= dataBufferIn(4068) when (flag_long='1') else '0';
	dataBufferOut(2173) <= dataBufferIn(4811) when (flag_long='1') else '0';
	dataBufferOut(2174) <= dataBufferIn(5554) when (flag_long='1') else '0';
	dataBufferOut(2175) <= dataBufferIn( 153) when (flag_long='1') else '0';
	dataBufferOut(2176) <= dataBufferIn( 896) when (flag_long='1') else '0';
	dataBufferOut(2177) <= dataBufferIn(1639) when (flag_long='1') else '0';
	dataBufferOut(2178) <= dataBufferIn(2382) when (flag_long='1') else '0';
	dataBufferOut(2179) <= dataBufferIn(3125) when (flag_long='1') else '0';
	dataBufferOut(2180) <= dataBufferIn(3868) when (flag_long='1') else '0';
	dataBufferOut(2181) <= dataBufferIn(4611) when (flag_long='1') else '0';
	dataBufferOut(2182) <= dataBufferIn(5354) when (flag_long='1') else '0';
	dataBufferOut(2183) <= dataBufferIn(6097) when (flag_long='1') else '0';
	dataBufferOut(2184) <= dataBufferIn( 696) when (flag_long='1') else '0';
	dataBufferOut(2185) <= dataBufferIn(1439) when (flag_long='1') else '0';
	dataBufferOut(2186) <= dataBufferIn(2182) when (flag_long='1') else '0';
	dataBufferOut(2187) <= dataBufferIn(2925) when (flag_long='1') else '0';
	dataBufferOut(2188) <= dataBufferIn(3668) when (flag_long='1') else '0';
	dataBufferOut(2189) <= dataBufferIn(4411) when (flag_long='1') else '0';
	dataBufferOut(2190) <= dataBufferIn(5154) when (flag_long='1') else '0';
	dataBufferOut(2191) <= dataBufferIn(5897) when (flag_long='1') else '0';
	dataBufferOut(2192) <= dataBufferIn( 496) when (flag_long='1') else '0';
	dataBufferOut(2193) <= dataBufferIn(1239) when (flag_long='1') else '0';
	dataBufferOut(2194) <= dataBufferIn(1982) when (flag_long='1') else '0';
	dataBufferOut(2195) <= dataBufferIn(2725) when (flag_long='1') else '0';
	dataBufferOut(2196) <= dataBufferIn(3468) when (flag_long='1') else '0';
	dataBufferOut(2197) <= dataBufferIn(4211) when (flag_long='1') else '0';
	dataBufferOut(2198) <= dataBufferIn(4954) when (flag_long='1') else '0';
	dataBufferOut(2199) <= dataBufferIn(5697) when (flag_long='1') else '0';
	dataBufferOut(2200) <= dataBufferIn( 296) when (flag_long='1') else '0';
	dataBufferOut(2201) <= dataBufferIn(1039) when (flag_long='1') else '0';
	dataBufferOut(2202) <= dataBufferIn(1782) when (flag_long='1') else '0';
	dataBufferOut(2203) <= dataBufferIn(2525) when (flag_long='1') else '0';
	dataBufferOut(2204) <= dataBufferIn(3268) when (flag_long='1') else '0';
	dataBufferOut(2205) <= dataBufferIn(4011) when (flag_long='1') else '0';
	dataBufferOut(2206) <= dataBufferIn(4754) when (flag_long='1') else '0';
	dataBufferOut(2207) <= dataBufferIn(5497) when (flag_long='1') else '0';
	dataBufferOut(2208) <= dataBufferIn(  96) when (flag_long='1') else '0';
	dataBufferOut(2209) <= dataBufferIn( 839) when (flag_long='1') else '0';
	dataBufferOut(2210) <= dataBufferIn(1582) when (flag_long='1') else '0';
	dataBufferOut(2211) <= dataBufferIn(2325) when (flag_long='1') else '0';
	dataBufferOut(2212) <= dataBufferIn(3068) when (flag_long='1') else '0';
	dataBufferOut(2213) <= dataBufferIn(3811) when (flag_long='1') else '0';
	dataBufferOut(2214) <= dataBufferIn(4554) when (flag_long='1') else '0';
	dataBufferOut(2215) <= dataBufferIn(5297) when (flag_long='1') else '0';
	dataBufferOut(2216) <= dataBufferIn(6040) when (flag_long='1') else '0';
	dataBufferOut(2217) <= dataBufferIn( 639) when (flag_long='1') else '0';
	dataBufferOut(2218) <= dataBufferIn(1382) when (flag_long='1') else '0';
	dataBufferOut(2219) <= dataBufferIn(2125) when (flag_long='1') else '0';
	dataBufferOut(2220) <= dataBufferIn(2868) when (flag_long='1') else '0';
	dataBufferOut(2221) <= dataBufferIn(3611) when (flag_long='1') else '0';
	dataBufferOut(2222) <= dataBufferIn(4354) when (flag_long='1') else '0';
	dataBufferOut(2223) <= dataBufferIn(5097) when (flag_long='1') else '0';
	dataBufferOut(2224) <= dataBufferIn(5840) when (flag_long='1') else '0';
	dataBufferOut(2225) <= dataBufferIn( 439) when (flag_long='1') else '0';
	dataBufferOut(2226) <= dataBufferIn(1182) when (flag_long='1') else '0';
	dataBufferOut(2227) <= dataBufferIn(1925) when (flag_long='1') else '0';
	dataBufferOut(2228) <= dataBufferIn(2668) when (flag_long='1') else '0';
	dataBufferOut(2229) <= dataBufferIn(3411) when (flag_long='1') else '0';
	dataBufferOut(2230) <= dataBufferIn(4154) when (flag_long='1') else '0';
	dataBufferOut(2231) <= dataBufferIn(4897) when (flag_long='1') else '0';
	dataBufferOut(2232) <= dataBufferIn(5640) when (flag_long='1') else '0';
	dataBufferOut(2233) <= dataBufferIn( 239) when (flag_long='1') else '0';
	dataBufferOut(2234) <= dataBufferIn( 982) when (flag_long='1') else '0';
	dataBufferOut(2235) <= dataBufferIn(1725) when (flag_long='1') else '0';
	dataBufferOut(2236) <= dataBufferIn(2468) when (flag_long='1') else '0';
	dataBufferOut(2237) <= dataBufferIn(3211) when (flag_long='1') else '0';
	dataBufferOut(2238) <= dataBufferIn(3954) when (flag_long='1') else '0';
	dataBufferOut(2239) <= dataBufferIn(4697) when (flag_long='1') else '0';
	dataBufferOut(2240) <= dataBufferIn(5440) when (flag_long='1') else '0';
	dataBufferOut(2241) <= dataBufferIn(  39) when (flag_long='1') else '0';
	dataBufferOut(2242) <= dataBufferIn( 782) when (flag_long='1') else '0';
	dataBufferOut(2243) <= dataBufferIn(1525) when (flag_long='1') else '0';
	dataBufferOut(2244) <= dataBufferIn(2268) when (flag_long='1') else '0';
	dataBufferOut(2245) <= dataBufferIn(3011) when (flag_long='1') else '0';
	dataBufferOut(2246) <= dataBufferIn(3754) when (flag_long='1') else '0';
	dataBufferOut(2247) <= dataBufferIn(4497) when (flag_long='1') else '0';
	dataBufferOut(2248) <= dataBufferIn(5240) when (flag_long='1') else '0';
	dataBufferOut(2249) <= dataBufferIn(5983) when (flag_long='1') else '0';
	dataBufferOut(2250) <= dataBufferIn( 582) when (flag_long='1') else '0';
	dataBufferOut(2251) <= dataBufferIn(1325) when (flag_long='1') else '0';
	dataBufferOut(2252) <= dataBufferIn(2068) when (flag_long='1') else '0';
	dataBufferOut(2253) <= dataBufferIn(2811) when (flag_long='1') else '0';
	dataBufferOut(2254) <= dataBufferIn(3554) when (flag_long='1') else '0';
	dataBufferOut(2255) <= dataBufferIn(4297) when (flag_long='1') else '0';
	dataBufferOut(2256) <= dataBufferIn(5040) when (flag_long='1') else '0';
	dataBufferOut(2257) <= dataBufferIn(5783) when (flag_long='1') else '0';
	dataBufferOut(2258) <= dataBufferIn( 382) when (flag_long='1') else '0';
	dataBufferOut(2259) <= dataBufferIn(1125) when (flag_long='1') else '0';
	dataBufferOut(2260) <= dataBufferIn(1868) when (flag_long='1') else '0';
	dataBufferOut(2261) <= dataBufferIn(2611) when (flag_long='1') else '0';
	dataBufferOut(2262) <= dataBufferIn(3354) when (flag_long='1') else '0';
	dataBufferOut(2263) <= dataBufferIn(4097) when (flag_long='1') else '0';
	dataBufferOut(2264) <= dataBufferIn(4840) when (flag_long='1') else '0';
	dataBufferOut(2265) <= dataBufferIn(5583) when (flag_long='1') else '0';
	dataBufferOut(2266) <= dataBufferIn( 182) when (flag_long='1') else '0';
	dataBufferOut(2267) <= dataBufferIn( 925) when (flag_long='1') else '0';
	dataBufferOut(2268) <= dataBufferIn(1668) when (flag_long='1') else '0';
	dataBufferOut(2269) <= dataBufferIn(2411) when (flag_long='1') else '0';
	dataBufferOut(2270) <= dataBufferIn(3154) when (flag_long='1') else '0';
	dataBufferOut(2271) <= dataBufferIn(3897) when (flag_long='1') else '0';
	dataBufferOut(2272) <= dataBufferIn(4640) when (flag_long='1') else '0';
	dataBufferOut(2273) <= dataBufferIn(5383) when (flag_long='1') else '0';
	dataBufferOut(2274) <= dataBufferIn(6126) when (flag_long='1') else '0';
	dataBufferOut(2275) <= dataBufferIn( 725) when (flag_long='1') else '0';
	dataBufferOut(2276) <= dataBufferIn(1468) when (flag_long='1') else '0';
	dataBufferOut(2277) <= dataBufferIn(2211) when (flag_long='1') else '0';
	dataBufferOut(2278) <= dataBufferIn(2954) when (flag_long='1') else '0';
	dataBufferOut(2279) <= dataBufferIn(3697) when (flag_long='1') else '0';
	dataBufferOut(2280) <= dataBufferIn(4440) when (flag_long='1') else '0';
	dataBufferOut(2281) <= dataBufferIn(5183) when (flag_long='1') else '0';
	dataBufferOut(2282) <= dataBufferIn(5926) when (flag_long='1') else '0';
	dataBufferOut(2283) <= dataBufferIn( 525) when (flag_long='1') else '0';
	dataBufferOut(2284) <= dataBufferIn(1268) when (flag_long='1') else '0';
	dataBufferOut(2285) <= dataBufferIn(2011) when (flag_long='1') else '0';
	dataBufferOut(2286) <= dataBufferIn(2754) when (flag_long='1') else '0';
	dataBufferOut(2287) <= dataBufferIn(3497) when (flag_long='1') else '0';
	dataBufferOut(2288) <= dataBufferIn(4240) when (flag_long='1') else '0';
	dataBufferOut(2289) <= dataBufferIn(4983) when (flag_long='1') else '0';
	dataBufferOut(2290) <= dataBufferIn(5726) when (flag_long='1') else '0';
	dataBufferOut(2291) <= dataBufferIn( 325) when (flag_long='1') else '0';
	dataBufferOut(2292) <= dataBufferIn(1068) when (flag_long='1') else '0';
	dataBufferOut(2293) <= dataBufferIn(1811) when (flag_long='1') else '0';
	dataBufferOut(2294) <= dataBufferIn(2554) when (flag_long='1') else '0';
	dataBufferOut(2295) <= dataBufferIn(3297) when (flag_long='1') else '0';
	dataBufferOut(2296) <= dataBufferIn(4040) when (flag_long='1') else '0';
	dataBufferOut(2297) <= dataBufferIn(4783) when (flag_long='1') else '0';
	dataBufferOut(2298) <= dataBufferIn(5526) when (flag_long='1') else '0';
	dataBufferOut(2299) <= dataBufferIn( 125) when (flag_long='1') else '0';
	dataBufferOut(2300) <= dataBufferIn( 868) when (flag_long='1') else '0';
	dataBufferOut(2301) <= dataBufferIn(1611) when (flag_long='1') else '0';
	dataBufferOut(2302) <= dataBufferIn(2354) when (flag_long='1') else '0';
	dataBufferOut(2303) <= dataBufferIn(3097) when (flag_long='1') else '0';
	dataBufferOut(2304) <= dataBufferIn(3840) when (flag_long='1') else '0';
	dataBufferOut(2305) <= dataBufferIn(4583) when (flag_long='1') else '0';
	dataBufferOut(2306) <= dataBufferIn(5326) when (flag_long='1') else '0';
	dataBufferOut(2307) <= dataBufferIn(6069) when (flag_long='1') else '0';
	dataBufferOut(2308) <= dataBufferIn( 668) when (flag_long='1') else '0';
	dataBufferOut(2309) <= dataBufferIn(1411) when (flag_long='1') else '0';
	dataBufferOut(2310) <= dataBufferIn(2154) when (flag_long='1') else '0';
	dataBufferOut(2311) <= dataBufferIn(2897) when (flag_long='1') else '0';
	dataBufferOut(2312) <= dataBufferIn(3640) when (flag_long='1') else '0';
	dataBufferOut(2313) <= dataBufferIn(4383) when (flag_long='1') else '0';
	dataBufferOut(2314) <= dataBufferIn(5126) when (flag_long='1') else '0';
	dataBufferOut(2315) <= dataBufferIn(5869) when (flag_long='1') else '0';
	dataBufferOut(2316) <= dataBufferIn( 468) when (flag_long='1') else '0';
	dataBufferOut(2317) <= dataBufferIn(1211) when (flag_long='1') else '0';
	dataBufferOut(2318) <= dataBufferIn(1954) when (flag_long='1') else '0';
	dataBufferOut(2319) <= dataBufferIn(2697) when (flag_long='1') else '0';
	dataBufferOut(2320) <= dataBufferIn(3440) when (flag_long='1') else '0';
	dataBufferOut(2321) <= dataBufferIn(4183) when (flag_long='1') else '0';
	dataBufferOut(2322) <= dataBufferIn(4926) when (flag_long='1') else '0';
	dataBufferOut(2323) <= dataBufferIn(5669) when (flag_long='1') else '0';
	dataBufferOut(2324) <= dataBufferIn( 268) when (flag_long='1') else '0';
	dataBufferOut(2325) <= dataBufferIn(1011) when (flag_long='1') else '0';
	dataBufferOut(2326) <= dataBufferIn(1754) when (flag_long='1') else '0';
	dataBufferOut(2327) <= dataBufferIn(2497) when (flag_long='1') else '0';
	dataBufferOut(2328) <= dataBufferIn(3240) when (flag_long='1') else '0';
	dataBufferOut(2329) <= dataBufferIn(3983) when (flag_long='1') else '0';
	dataBufferOut(2330) <= dataBufferIn(4726) when (flag_long='1') else '0';
	dataBufferOut(2331) <= dataBufferIn(5469) when (flag_long='1') else '0';
	dataBufferOut(2332) <= dataBufferIn(  68) when (flag_long='1') else '0';
	dataBufferOut(2333) <= dataBufferIn( 811) when (flag_long='1') else '0';
	dataBufferOut(2334) <= dataBufferIn(1554) when (flag_long='1') else '0';
	dataBufferOut(2335) <= dataBufferIn(2297) when (flag_long='1') else '0';
	dataBufferOut(2336) <= dataBufferIn(3040) when (flag_long='1') else '0';
	dataBufferOut(2337) <= dataBufferIn(3783) when (flag_long='1') else '0';
	dataBufferOut(2338) <= dataBufferIn(4526) when (flag_long='1') else '0';
	dataBufferOut(2339) <= dataBufferIn(5269) when (flag_long='1') else '0';
	dataBufferOut(2340) <= dataBufferIn(6012) when (flag_long='1') else '0';
	dataBufferOut(2341) <= dataBufferIn( 611) when (flag_long='1') else '0';
	dataBufferOut(2342) <= dataBufferIn(1354) when (flag_long='1') else '0';
	dataBufferOut(2343) <= dataBufferIn(2097) when (flag_long='1') else '0';
	dataBufferOut(2344) <= dataBufferIn(2840) when (flag_long='1') else '0';
	dataBufferOut(2345) <= dataBufferIn(3583) when (flag_long='1') else '0';
	dataBufferOut(2346) <= dataBufferIn(4326) when (flag_long='1') else '0';
	dataBufferOut(2347) <= dataBufferIn(5069) when (flag_long='1') else '0';
	dataBufferOut(2348) <= dataBufferIn(5812) when (flag_long='1') else '0';
	dataBufferOut(2349) <= dataBufferIn( 411) when (flag_long='1') else '0';
	dataBufferOut(2350) <= dataBufferIn(1154) when (flag_long='1') else '0';
	dataBufferOut(2351) <= dataBufferIn(1897) when (flag_long='1') else '0';
	dataBufferOut(2352) <= dataBufferIn(2640) when (flag_long='1') else '0';
	dataBufferOut(2353) <= dataBufferIn(3383) when (flag_long='1') else '0';
	dataBufferOut(2354) <= dataBufferIn(4126) when (flag_long='1') else '0';
	dataBufferOut(2355) <= dataBufferIn(4869) when (flag_long='1') else '0';
	dataBufferOut(2356) <= dataBufferIn(5612) when (flag_long='1') else '0';
	dataBufferOut(2357) <= dataBufferIn( 211) when (flag_long='1') else '0';
	dataBufferOut(2358) <= dataBufferIn( 954) when (flag_long='1') else '0';
	dataBufferOut(2359) <= dataBufferIn(1697) when (flag_long='1') else '0';
	dataBufferOut(2360) <= dataBufferIn(2440) when (flag_long='1') else '0';
	dataBufferOut(2361) <= dataBufferIn(3183) when (flag_long='1') else '0';
	dataBufferOut(2362) <= dataBufferIn(3926) when (flag_long='1') else '0';
	dataBufferOut(2363) <= dataBufferIn(4669) when (flag_long='1') else '0';
	dataBufferOut(2364) <= dataBufferIn(5412) when (flag_long='1') else '0';
	dataBufferOut(2365) <= dataBufferIn(  11) when (flag_long='1') else '0';
	dataBufferOut(2366) <= dataBufferIn( 754) when (flag_long='1') else '0';
	dataBufferOut(2367) <= dataBufferIn(1497) when (flag_long='1') else '0';
	dataBufferOut(2368) <= dataBufferIn(2240) when (flag_long='1') else '0';
	dataBufferOut(2369) <= dataBufferIn(2983) when (flag_long='1') else '0';
	dataBufferOut(2370) <= dataBufferIn(3726) when (flag_long='1') else '0';
	dataBufferOut(2371) <= dataBufferIn(4469) when (flag_long='1') else '0';
	dataBufferOut(2372) <= dataBufferIn(5212) when (flag_long='1') else '0';
	dataBufferOut(2373) <= dataBufferIn(5955) when (flag_long='1') else '0';
	dataBufferOut(2374) <= dataBufferIn( 554) when (flag_long='1') else '0';
	dataBufferOut(2375) <= dataBufferIn(1297) when (flag_long='1') else '0';
	dataBufferOut(2376) <= dataBufferIn(2040) when (flag_long='1') else '0';
	dataBufferOut(2377) <= dataBufferIn(2783) when (flag_long='1') else '0';
	dataBufferOut(2378) <= dataBufferIn(3526) when (flag_long='1') else '0';
	dataBufferOut(2379) <= dataBufferIn(4269) when (flag_long='1') else '0';
	dataBufferOut(2380) <= dataBufferIn(5012) when (flag_long='1') else '0';
	dataBufferOut(2381) <= dataBufferIn(5755) when (flag_long='1') else '0';
	dataBufferOut(2382) <= dataBufferIn( 354) when (flag_long='1') else '0';
	dataBufferOut(2383) <= dataBufferIn(1097) when (flag_long='1') else '0';
	dataBufferOut(2384) <= dataBufferIn(1840) when (flag_long='1') else '0';
	dataBufferOut(2385) <= dataBufferIn(2583) when (flag_long='1') else '0';
	dataBufferOut(2386) <= dataBufferIn(3326) when (flag_long='1') else '0';
	dataBufferOut(2387) <= dataBufferIn(4069) when (flag_long='1') else '0';
	dataBufferOut(2388) <= dataBufferIn(4812) when (flag_long='1') else '0';
	dataBufferOut(2389) <= dataBufferIn(5555) when (flag_long='1') else '0';
	dataBufferOut(2390) <= dataBufferIn( 154) when (flag_long='1') else '0';
	dataBufferOut(2391) <= dataBufferIn( 897) when (flag_long='1') else '0';
	dataBufferOut(2392) <= dataBufferIn(1640) when (flag_long='1') else '0';
	dataBufferOut(2393) <= dataBufferIn(2383) when (flag_long='1') else '0';
	dataBufferOut(2394) <= dataBufferIn(3126) when (flag_long='1') else '0';
	dataBufferOut(2395) <= dataBufferIn(3869) when (flag_long='1') else '0';
	dataBufferOut(2396) <= dataBufferIn(4612) when (flag_long='1') else '0';
	dataBufferOut(2397) <= dataBufferIn(5355) when (flag_long='1') else '0';
	dataBufferOut(2398) <= dataBufferIn(6098) when (flag_long='1') else '0';
	dataBufferOut(2399) <= dataBufferIn( 697) when (flag_long='1') else '0';
	dataBufferOut(2400) <= dataBufferIn(1440) when (flag_long='1') else '0';
	dataBufferOut(2401) <= dataBufferIn(2183) when (flag_long='1') else '0';
	dataBufferOut(2402) <= dataBufferIn(2926) when (flag_long='1') else '0';
	dataBufferOut(2403) <= dataBufferIn(3669) when (flag_long='1') else '0';
	dataBufferOut(2404) <= dataBufferIn(4412) when (flag_long='1') else '0';
	dataBufferOut(2405) <= dataBufferIn(5155) when (flag_long='1') else '0';
	dataBufferOut(2406) <= dataBufferIn(5898) when (flag_long='1') else '0';
	dataBufferOut(2407) <= dataBufferIn( 497) when (flag_long='1') else '0';
	dataBufferOut(2408) <= dataBufferIn(1240) when (flag_long='1') else '0';
	dataBufferOut(2409) <= dataBufferIn(1983) when (flag_long='1') else '0';
	dataBufferOut(2410) <= dataBufferIn(2726) when (flag_long='1') else '0';
	dataBufferOut(2411) <= dataBufferIn(3469) when (flag_long='1') else '0';
	dataBufferOut(2412) <= dataBufferIn(4212) when (flag_long='1') else '0';
	dataBufferOut(2413) <= dataBufferIn(4955) when (flag_long='1') else '0';
	dataBufferOut(2414) <= dataBufferIn(5698) when (flag_long='1') else '0';
	dataBufferOut(2415) <= dataBufferIn( 297) when (flag_long='1') else '0';
	dataBufferOut(2416) <= dataBufferIn(1040) when (flag_long='1') else '0';
	dataBufferOut(2417) <= dataBufferIn(1783) when (flag_long='1') else '0';
	dataBufferOut(2418) <= dataBufferIn(2526) when (flag_long='1') else '0';
	dataBufferOut(2419) <= dataBufferIn(3269) when (flag_long='1') else '0';
	dataBufferOut(2420) <= dataBufferIn(4012) when (flag_long='1') else '0';
	dataBufferOut(2421) <= dataBufferIn(4755) when (flag_long='1') else '0';
	dataBufferOut(2422) <= dataBufferIn(5498) when (flag_long='1') else '0';
	dataBufferOut(2423) <= dataBufferIn(  97) when (flag_long='1') else '0';
	dataBufferOut(2424) <= dataBufferIn( 840) when (flag_long='1') else '0';
	dataBufferOut(2425) <= dataBufferIn(1583) when (flag_long='1') else '0';
	dataBufferOut(2426) <= dataBufferIn(2326) when (flag_long='1') else '0';
	dataBufferOut(2427) <= dataBufferIn(3069) when (flag_long='1') else '0';
	dataBufferOut(2428) <= dataBufferIn(3812) when (flag_long='1') else '0';
	dataBufferOut(2429) <= dataBufferIn(4555) when (flag_long='1') else '0';
	dataBufferOut(2430) <= dataBufferIn(5298) when (flag_long='1') else '0';
	dataBufferOut(2431) <= dataBufferIn(6041) when (flag_long='1') else '0';
	dataBufferOut(2432) <= dataBufferIn( 640) when (flag_long='1') else '0';
	dataBufferOut(2433) <= dataBufferIn(1383) when (flag_long='1') else '0';
	dataBufferOut(2434) <= dataBufferIn(2126) when (flag_long='1') else '0';
	dataBufferOut(2435) <= dataBufferIn(2869) when (flag_long='1') else '0';
	dataBufferOut(2436) <= dataBufferIn(3612) when (flag_long='1') else '0';
	dataBufferOut(2437) <= dataBufferIn(4355) when (flag_long='1') else '0';
	dataBufferOut(2438) <= dataBufferIn(5098) when (flag_long='1') else '0';
	dataBufferOut(2439) <= dataBufferIn(5841) when (flag_long='1') else '0';
	dataBufferOut(2440) <= dataBufferIn( 440) when (flag_long='1') else '0';
	dataBufferOut(2441) <= dataBufferIn(1183) when (flag_long='1') else '0';
	dataBufferOut(2442) <= dataBufferIn(1926) when (flag_long='1') else '0';
	dataBufferOut(2443) <= dataBufferIn(2669) when (flag_long='1') else '0';
	dataBufferOut(2444) <= dataBufferIn(3412) when (flag_long='1') else '0';
	dataBufferOut(2445) <= dataBufferIn(4155) when (flag_long='1') else '0';
	dataBufferOut(2446) <= dataBufferIn(4898) when (flag_long='1') else '0';
	dataBufferOut(2447) <= dataBufferIn(5641) when (flag_long='1') else '0';
	dataBufferOut(2448) <= dataBufferIn( 240) when (flag_long='1') else '0';
	dataBufferOut(2449) <= dataBufferIn( 983) when (flag_long='1') else '0';
	dataBufferOut(2450) <= dataBufferIn(1726) when (flag_long='1') else '0';
	dataBufferOut(2451) <= dataBufferIn(2469) when (flag_long='1') else '0';
	dataBufferOut(2452) <= dataBufferIn(3212) when (flag_long='1') else '0';
	dataBufferOut(2453) <= dataBufferIn(3955) when (flag_long='1') else '0';
	dataBufferOut(2454) <= dataBufferIn(4698) when (flag_long='1') else '0';
	dataBufferOut(2455) <= dataBufferIn(5441) when (flag_long='1') else '0';
	dataBufferOut(2456) <= dataBufferIn(  40) when (flag_long='1') else '0';
	dataBufferOut(2457) <= dataBufferIn( 783) when (flag_long='1') else '0';
	dataBufferOut(2458) <= dataBufferIn(1526) when (flag_long='1') else '0';
	dataBufferOut(2459) <= dataBufferIn(2269) when (flag_long='1') else '0';
	dataBufferOut(2460) <= dataBufferIn(3012) when (flag_long='1') else '0';
	dataBufferOut(2461) <= dataBufferIn(3755) when (flag_long='1') else '0';
	dataBufferOut(2462) <= dataBufferIn(4498) when (flag_long='1') else '0';
	dataBufferOut(2463) <= dataBufferIn(5241) when (flag_long='1') else '0';
	dataBufferOut(2464) <= dataBufferIn(5984) when (flag_long='1') else '0';
	dataBufferOut(2465) <= dataBufferIn( 583) when (flag_long='1') else '0';
	dataBufferOut(2466) <= dataBufferIn(1326) when (flag_long='1') else '0';
	dataBufferOut(2467) <= dataBufferIn(2069) when (flag_long='1') else '0';
	dataBufferOut(2468) <= dataBufferIn(2812) when (flag_long='1') else '0';
	dataBufferOut(2469) <= dataBufferIn(3555) when (flag_long='1') else '0';
	dataBufferOut(2470) <= dataBufferIn(4298) when (flag_long='1') else '0';
	dataBufferOut(2471) <= dataBufferIn(5041) when (flag_long='1') else '0';
	dataBufferOut(2472) <= dataBufferIn(5784) when (flag_long='1') else '0';
	dataBufferOut(2473) <= dataBufferIn( 383) when (flag_long='1') else '0';
	dataBufferOut(2474) <= dataBufferIn(1126) when (flag_long='1') else '0';
	dataBufferOut(2475) <= dataBufferIn(1869) when (flag_long='1') else '0';
	dataBufferOut(2476) <= dataBufferIn(2612) when (flag_long='1') else '0';
	dataBufferOut(2477) <= dataBufferIn(3355) when (flag_long='1') else '0';
	dataBufferOut(2478) <= dataBufferIn(4098) when (flag_long='1') else '0';
	dataBufferOut(2479) <= dataBufferIn(4841) when (flag_long='1') else '0';
	dataBufferOut(2480) <= dataBufferIn(5584) when (flag_long='1') else '0';
	dataBufferOut(2481) <= dataBufferIn( 183) when (flag_long='1') else '0';
	dataBufferOut(2482) <= dataBufferIn( 926) when (flag_long='1') else '0';
	dataBufferOut(2483) <= dataBufferIn(1669) when (flag_long='1') else '0';
	dataBufferOut(2484) <= dataBufferIn(2412) when (flag_long='1') else '0';
	dataBufferOut(2485) <= dataBufferIn(3155) when (flag_long='1') else '0';
	dataBufferOut(2486) <= dataBufferIn(3898) when (flag_long='1') else '0';
	dataBufferOut(2487) <= dataBufferIn(4641) when (flag_long='1') else '0';
	dataBufferOut(2488) <= dataBufferIn(5384) when (flag_long='1') else '0';
	dataBufferOut(2489) <= dataBufferIn(6127) when (flag_long='1') else '0';
	dataBufferOut(2490) <= dataBufferIn( 726) when (flag_long='1') else '0';
	dataBufferOut(2491) <= dataBufferIn(1469) when (flag_long='1') else '0';
	dataBufferOut(2492) <= dataBufferIn(2212) when (flag_long='1') else '0';
	dataBufferOut(2493) <= dataBufferIn(2955) when (flag_long='1') else '0';
	dataBufferOut(2494) <= dataBufferIn(3698) when (flag_long='1') else '0';
	dataBufferOut(2495) <= dataBufferIn(4441) when (flag_long='1') else '0';
	dataBufferOut(2496) <= dataBufferIn(5184) when (flag_long='1') else '0';
	dataBufferOut(2497) <= dataBufferIn(5927) when (flag_long='1') else '0';
	dataBufferOut(2498) <= dataBufferIn( 526) when (flag_long='1') else '0';
	dataBufferOut(2499) <= dataBufferIn(1269) when (flag_long='1') else '0';
	dataBufferOut(2500) <= dataBufferIn(2012) when (flag_long='1') else '0';
	dataBufferOut(2501) <= dataBufferIn(2755) when (flag_long='1') else '0';
	dataBufferOut(2502) <= dataBufferIn(3498) when (flag_long='1') else '0';
	dataBufferOut(2503) <= dataBufferIn(4241) when (flag_long='1') else '0';
	dataBufferOut(2504) <= dataBufferIn(4984) when (flag_long='1') else '0';
	dataBufferOut(2505) <= dataBufferIn(5727) when (flag_long='1') else '0';
	dataBufferOut(2506) <= dataBufferIn( 326) when (flag_long='1') else '0';
	dataBufferOut(2507) <= dataBufferIn(1069) when (flag_long='1') else '0';
	dataBufferOut(2508) <= dataBufferIn(1812) when (flag_long='1') else '0';
	dataBufferOut(2509) <= dataBufferIn(2555) when (flag_long='1') else '0';
	dataBufferOut(2510) <= dataBufferIn(3298) when (flag_long='1') else '0';
	dataBufferOut(2511) <= dataBufferIn(4041) when (flag_long='1') else '0';
	dataBufferOut(2512) <= dataBufferIn(4784) when (flag_long='1') else '0';
	dataBufferOut(2513) <= dataBufferIn(5527) when (flag_long='1') else '0';
	dataBufferOut(2514) <= dataBufferIn( 126) when (flag_long='1') else '0';
	dataBufferOut(2515) <= dataBufferIn( 869) when (flag_long='1') else '0';
	dataBufferOut(2516) <= dataBufferIn(1612) when (flag_long='1') else '0';
	dataBufferOut(2517) <= dataBufferIn(2355) when (flag_long='1') else '0';
	dataBufferOut(2518) <= dataBufferIn(3098) when (flag_long='1') else '0';
	dataBufferOut(2519) <= dataBufferIn(3841) when (flag_long='1') else '0';
	dataBufferOut(2520) <= dataBufferIn(4584) when (flag_long='1') else '0';
	dataBufferOut(2521) <= dataBufferIn(5327) when (flag_long='1') else '0';
	dataBufferOut(2522) <= dataBufferIn(6070) when (flag_long='1') else '0';
	dataBufferOut(2523) <= dataBufferIn( 669) when (flag_long='1') else '0';
	dataBufferOut(2524) <= dataBufferIn(1412) when (flag_long='1') else '0';
	dataBufferOut(2525) <= dataBufferIn(2155) when (flag_long='1') else '0';
	dataBufferOut(2526) <= dataBufferIn(2898) when (flag_long='1') else '0';
	dataBufferOut(2527) <= dataBufferIn(3641) when (flag_long='1') else '0';
	dataBufferOut(2528) <= dataBufferIn(4384) when (flag_long='1') else '0';
	dataBufferOut(2529) <= dataBufferIn(5127) when (flag_long='1') else '0';
	dataBufferOut(2530) <= dataBufferIn(5870) when (flag_long='1') else '0';
	dataBufferOut(2531) <= dataBufferIn( 469) when (flag_long='1') else '0';
	dataBufferOut(2532) <= dataBufferIn(1212) when (flag_long='1') else '0';
	dataBufferOut(2533) <= dataBufferIn(1955) when (flag_long='1') else '0';
	dataBufferOut(2534) <= dataBufferIn(2698) when (flag_long='1') else '0';
	dataBufferOut(2535) <= dataBufferIn(3441) when (flag_long='1') else '0';
	dataBufferOut(2536) <= dataBufferIn(4184) when (flag_long='1') else '0';
	dataBufferOut(2537) <= dataBufferIn(4927) when (flag_long='1') else '0';
	dataBufferOut(2538) <= dataBufferIn(5670) when (flag_long='1') else '0';
	dataBufferOut(2539) <= dataBufferIn( 269) when (flag_long='1') else '0';
	dataBufferOut(2540) <= dataBufferIn(1012) when (flag_long='1') else '0';
	dataBufferOut(2541) <= dataBufferIn(1755) when (flag_long='1') else '0';
	dataBufferOut(2542) <= dataBufferIn(2498) when (flag_long='1') else '0';
	dataBufferOut(2543) <= dataBufferIn(3241) when (flag_long='1') else '0';
	dataBufferOut(2544) <= dataBufferIn(3984) when (flag_long='1') else '0';
	dataBufferOut(2545) <= dataBufferIn(4727) when (flag_long='1') else '0';
	dataBufferOut(2546) <= dataBufferIn(5470) when (flag_long='1') else '0';
	dataBufferOut(2547) <= dataBufferIn(  69) when (flag_long='1') else '0';
	dataBufferOut(2548) <= dataBufferIn( 812) when (flag_long='1') else '0';
	dataBufferOut(2549) <= dataBufferIn(1555) when (flag_long='1') else '0';
	dataBufferOut(2550) <= dataBufferIn(2298) when (flag_long='1') else '0';
	dataBufferOut(2551) <= dataBufferIn(3041) when (flag_long='1') else '0';
	dataBufferOut(2552) <= dataBufferIn(3784) when (flag_long='1') else '0';
	dataBufferOut(2553) <= dataBufferIn(4527) when (flag_long='1') else '0';
	dataBufferOut(2554) <= dataBufferIn(5270) when (flag_long='1') else '0';
	dataBufferOut(2555) <= dataBufferIn(6013) when (flag_long='1') else '0';
	dataBufferOut(2556) <= dataBufferIn( 612) when (flag_long='1') else '0';
	dataBufferOut(2557) <= dataBufferIn(1355) when (flag_long='1') else '0';
	dataBufferOut(2558) <= dataBufferIn(2098) when (flag_long='1') else '0';
	dataBufferOut(2559) <= dataBufferIn(2841) when (flag_long='1') else '0';
	dataBufferOut(2560) <= dataBufferIn(3584) when (flag_long='1') else '0';
	dataBufferOut(2561) <= dataBufferIn(4327) when (flag_long='1') else '0';
	dataBufferOut(2562) <= dataBufferIn(5070) when (flag_long='1') else '0';
	dataBufferOut(2563) <= dataBufferIn(5813) when (flag_long='1') else '0';
	dataBufferOut(2564) <= dataBufferIn( 412) when (flag_long='1') else '0';
	dataBufferOut(2565) <= dataBufferIn(1155) when (flag_long='1') else '0';
	dataBufferOut(2566) <= dataBufferIn(1898) when (flag_long='1') else '0';
	dataBufferOut(2567) <= dataBufferIn(2641) when (flag_long='1') else '0';
	dataBufferOut(2568) <= dataBufferIn(3384) when (flag_long='1') else '0';
	dataBufferOut(2569) <= dataBufferIn(4127) when (flag_long='1') else '0';
	dataBufferOut(2570) <= dataBufferIn(4870) when (flag_long='1') else '0';
	dataBufferOut(2571) <= dataBufferIn(5613) when (flag_long='1') else '0';
	dataBufferOut(2572) <= dataBufferIn( 212) when (flag_long='1') else '0';
	dataBufferOut(2573) <= dataBufferIn( 955) when (flag_long='1') else '0';
	dataBufferOut(2574) <= dataBufferIn(1698) when (flag_long='1') else '0';
	dataBufferOut(2575) <= dataBufferIn(2441) when (flag_long='1') else '0';
	dataBufferOut(2576) <= dataBufferIn(3184) when (flag_long='1') else '0';
	dataBufferOut(2577) <= dataBufferIn(3927) when (flag_long='1') else '0';
	dataBufferOut(2578) <= dataBufferIn(4670) when (flag_long='1') else '0';
	dataBufferOut(2579) <= dataBufferIn(5413) when (flag_long='1') else '0';
	dataBufferOut(2580) <= dataBufferIn(  12) when (flag_long='1') else '0';
	dataBufferOut(2581) <= dataBufferIn( 755) when (flag_long='1') else '0';
	dataBufferOut(2582) <= dataBufferIn(1498) when (flag_long='1') else '0';
	dataBufferOut(2583) <= dataBufferIn(2241) when (flag_long='1') else '0';
	dataBufferOut(2584) <= dataBufferIn(2984) when (flag_long='1') else '0';
	dataBufferOut(2585) <= dataBufferIn(3727) when (flag_long='1') else '0';
	dataBufferOut(2586) <= dataBufferIn(4470) when (flag_long='1') else '0';
	dataBufferOut(2587) <= dataBufferIn(5213) when (flag_long='1') else '0';
	dataBufferOut(2588) <= dataBufferIn(5956) when (flag_long='1') else '0';
	dataBufferOut(2589) <= dataBufferIn( 555) when (flag_long='1') else '0';
	dataBufferOut(2590) <= dataBufferIn(1298) when (flag_long='1') else '0';
	dataBufferOut(2591) <= dataBufferIn(2041) when (flag_long='1') else '0';
	dataBufferOut(2592) <= dataBufferIn(2784) when (flag_long='1') else '0';
	dataBufferOut(2593) <= dataBufferIn(3527) when (flag_long='1') else '0';
	dataBufferOut(2594) <= dataBufferIn(4270) when (flag_long='1') else '0';
	dataBufferOut(2595) <= dataBufferIn(5013) when (flag_long='1') else '0';
	dataBufferOut(2596) <= dataBufferIn(5756) when (flag_long='1') else '0';
	dataBufferOut(2597) <= dataBufferIn( 355) when (flag_long='1') else '0';
	dataBufferOut(2598) <= dataBufferIn(1098) when (flag_long='1') else '0';
	dataBufferOut(2599) <= dataBufferIn(1841) when (flag_long='1') else '0';
	dataBufferOut(2600) <= dataBufferIn(2584) when (flag_long='1') else '0';
	dataBufferOut(2601) <= dataBufferIn(3327) when (flag_long='1') else '0';
	dataBufferOut(2602) <= dataBufferIn(4070) when (flag_long='1') else '0';
	dataBufferOut(2603) <= dataBufferIn(4813) when (flag_long='1') else '0';
	dataBufferOut(2604) <= dataBufferIn(5556) when (flag_long='1') else '0';
	dataBufferOut(2605) <= dataBufferIn( 155) when (flag_long='1') else '0';
	dataBufferOut(2606) <= dataBufferIn( 898) when (flag_long='1') else '0';
	dataBufferOut(2607) <= dataBufferIn(1641) when (flag_long='1') else '0';
	dataBufferOut(2608) <= dataBufferIn(2384) when (flag_long='1') else '0';
	dataBufferOut(2609) <= dataBufferIn(3127) when (flag_long='1') else '0';
	dataBufferOut(2610) <= dataBufferIn(3870) when (flag_long='1') else '0';
	dataBufferOut(2611) <= dataBufferIn(4613) when (flag_long='1') else '0';
	dataBufferOut(2612) <= dataBufferIn(5356) when (flag_long='1') else '0';
	dataBufferOut(2613) <= dataBufferIn(6099) when (flag_long='1') else '0';
	dataBufferOut(2614) <= dataBufferIn( 698) when (flag_long='1') else '0';
	dataBufferOut(2615) <= dataBufferIn(1441) when (flag_long='1') else '0';
	dataBufferOut(2616) <= dataBufferIn(2184) when (flag_long='1') else '0';
	dataBufferOut(2617) <= dataBufferIn(2927) when (flag_long='1') else '0';
	dataBufferOut(2618) <= dataBufferIn(3670) when (flag_long='1') else '0';
	dataBufferOut(2619) <= dataBufferIn(4413) when (flag_long='1') else '0';
	dataBufferOut(2620) <= dataBufferIn(5156) when (flag_long='1') else '0';
	dataBufferOut(2621) <= dataBufferIn(5899) when (flag_long='1') else '0';
	dataBufferOut(2622) <= dataBufferIn( 498) when (flag_long='1') else '0';
	dataBufferOut(2623) <= dataBufferIn(1241) when (flag_long='1') else '0';
	dataBufferOut(2624) <= dataBufferIn(1984) when (flag_long='1') else '0';
	dataBufferOut(2625) <= dataBufferIn(2727) when (flag_long='1') else '0';
	dataBufferOut(2626) <= dataBufferIn(3470) when (flag_long='1') else '0';
	dataBufferOut(2627) <= dataBufferIn(4213) when (flag_long='1') else '0';
	dataBufferOut(2628) <= dataBufferIn(4956) when (flag_long='1') else '0';
	dataBufferOut(2629) <= dataBufferIn(5699) when (flag_long='1') else '0';
	dataBufferOut(2630) <= dataBufferIn( 298) when (flag_long='1') else '0';
	dataBufferOut(2631) <= dataBufferIn(1041) when (flag_long='1') else '0';
	dataBufferOut(2632) <= dataBufferIn(1784) when (flag_long='1') else '0';
	dataBufferOut(2633) <= dataBufferIn(2527) when (flag_long='1') else '0';
	dataBufferOut(2634) <= dataBufferIn(3270) when (flag_long='1') else '0';
	dataBufferOut(2635) <= dataBufferIn(4013) when (flag_long='1') else '0';
	dataBufferOut(2636) <= dataBufferIn(4756) when (flag_long='1') else '0';
	dataBufferOut(2637) <= dataBufferIn(5499) when (flag_long='1') else '0';
	dataBufferOut(2638) <= dataBufferIn(  98) when (flag_long='1') else '0';
	dataBufferOut(2639) <= dataBufferIn( 841) when (flag_long='1') else '0';
	dataBufferOut(2640) <= dataBufferIn(1584) when (flag_long='1') else '0';
	dataBufferOut(2641) <= dataBufferIn(2327) when (flag_long='1') else '0';
	dataBufferOut(2642) <= dataBufferIn(3070) when (flag_long='1') else '0';
	dataBufferOut(2643) <= dataBufferIn(3813) when (flag_long='1') else '0';
	dataBufferOut(2644) <= dataBufferIn(4556) when (flag_long='1') else '0';
	dataBufferOut(2645) <= dataBufferIn(5299) when (flag_long='1') else '0';
	dataBufferOut(2646) <= dataBufferIn(6042) when (flag_long='1') else '0';
	dataBufferOut(2647) <= dataBufferIn( 641) when (flag_long='1') else '0';
	dataBufferOut(2648) <= dataBufferIn(1384) when (flag_long='1') else '0';
	dataBufferOut(2649) <= dataBufferIn(2127) when (flag_long='1') else '0';
	dataBufferOut(2650) <= dataBufferIn(2870) when (flag_long='1') else '0';
	dataBufferOut(2651) <= dataBufferIn(3613) when (flag_long='1') else '0';
	dataBufferOut(2652) <= dataBufferIn(4356) when (flag_long='1') else '0';
	dataBufferOut(2653) <= dataBufferIn(5099) when (flag_long='1') else '0';
	dataBufferOut(2654) <= dataBufferIn(5842) when (flag_long='1') else '0';
	dataBufferOut(2655) <= dataBufferIn( 441) when (flag_long='1') else '0';
	dataBufferOut(2656) <= dataBufferIn(1184) when (flag_long='1') else '0';
	dataBufferOut(2657) <= dataBufferIn(1927) when (flag_long='1') else '0';
	dataBufferOut(2658) <= dataBufferIn(2670) when (flag_long='1') else '0';
	dataBufferOut(2659) <= dataBufferIn(3413) when (flag_long='1') else '0';
	dataBufferOut(2660) <= dataBufferIn(4156) when (flag_long='1') else '0';
	dataBufferOut(2661) <= dataBufferIn(4899) when (flag_long='1') else '0';
	dataBufferOut(2662) <= dataBufferIn(5642) when (flag_long='1') else '0';
	dataBufferOut(2663) <= dataBufferIn( 241) when (flag_long='1') else '0';
	dataBufferOut(2664) <= dataBufferIn( 984) when (flag_long='1') else '0';
	dataBufferOut(2665) <= dataBufferIn(1727) when (flag_long='1') else '0';
	dataBufferOut(2666) <= dataBufferIn(2470) when (flag_long='1') else '0';
	dataBufferOut(2667) <= dataBufferIn(3213) when (flag_long='1') else '0';
	dataBufferOut(2668) <= dataBufferIn(3956) when (flag_long='1') else '0';
	dataBufferOut(2669) <= dataBufferIn(4699) when (flag_long='1') else '0';
	dataBufferOut(2670) <= dataBufferIn(5442) when (flag_long='1') else '0';
	dataBufferOut(2671) <= dataBufferIn(  41) when (flag_long='1') else '0';
	dataBufferOut(2672) <= dataBufferIn( 784) when (flag_long='1') else '0';
	dataBufferOut(2673) <= dataBufferIn(1527) when (flag_long='1') else '0';
	dataBufferOut(2674) <= dataBufferIn(2270) when (flag_long='1') else '0';
	dataBufferOut(2675) <= dataBufferIn(3013) when (flag_long='1') else '0';
	dataBufferOut(2676) <= dataBufferIn(3756) when (flag_long='1') else '0';
	dataBufferOut(2677) <= dataBufferIn(4499) when (flag_long='1') else '0';
	dataBufferOut(2678) <= dataBufferIn(5242) when (flag_long='1') else '0';
	dataBufferOut(2679) <= dataBufferIn(5985) when (flag_long='1') else '0';
	dataBufferOut(2680) <= dataBufferIn( 584) when (flag_long='1') else '0';
	dataBufferOut(2681) <= dataBufferIn(1327) when (flag_long='1') else '0';
	dataBufferOut(2682) <= dataBufferIn(2070) when (flag_long='1') else '0';
	dataBufferOut(2683) <= dataBufferIn(2813) when (flag_long='1') else '0';
	dataBufferOut(2684) <= dataBufferIn(3556) when (flag_long='1') else '0';
	dataBufferOut(2685) <= dataBufferIn(4299) when (flag_long='1') else '0';
	dataBufferOut(2686) <= dataBufferIn(5042) when (flag_long='1') else '0';
	dataBufferOut(2687) <= dataBufferIn(5785) when (flag_long='1') else '0';
	dataBufferOut(2688) <= dataBufferIn( 384) when (flag_long='1') else '0';
	dataBufferOut(2689) <= dataBufferIn(1127) when (flag_long='1') else '0';
	dataBufferOut(2690) <= dataBufferIn(1870) when (flag_long='1') else '0';
	dataBufferOut(2691) <= dataBufferIn(2613) when (flag_long='1') else '0';
	dataBufferOut(2692) <= dataBufferIn(3356) when (flag_long='1') else '0';
	dataBufferOut(2693) <= dataBufferIn(4099) when (flag_long='1') else '0';
	dataBufferOut(2694) <= dataBufferIn(4842) when (flag_long='1') else '0';
	dataBufferOut(2695) <= dataBufferIn(5585) when (flag_long='1') else '0';
	dataBufferOut(2696) <= dataBufferIn( 184) when (flag_long='1') else '0';
	dataBufferOut(2697) <= dataBufferIn( 927) when (flag_long='1') else '0';
	dataBufferOut(2698) <= dataBufferIn(1670) when (flag_long='1') else '0';
	dataBufferOut(2699) <= dataBufferIn(2413) when (flag_long='1') else '0';
	dataBufferOut(2700) <= dataBufferIn(3156) when (flag_long='1') else '0';
	dataBufferOut(2701) <= dataBufferIn(3899) when (flag_long='1') else '0';
	dataBufferOut(2702) <= dataBufferIn(4642) when (flag_long='1') else '0';
	dataBufferOut(2703) <= dataBufferIn(5385) when (flag_long='1') else '0';
	dataBufferOut(2704) <= dataBufferIn(6128) when (flag_long='1') else '0';
	dataBufferOut(2705) <= dataBufferIn( 727) when (flag_long='1') else '0';
	dataBufferOut(2706) <= dataBufferIn(1470) when (flag_long='1') else '0';
	dataBufferOut(2707) <= dataBufferIn(2213) when (flag_long='1') else '0';
	dataBufferOut(2708) <= dataBufferIn(2956) when (flag_long='1') else '0';
	dataBufferOut(2709) <= dataBufferIn(3699) when (flag_long='1') else '0';
	dataBufferOut(2710) <= dataBufferIn(4442) when (flag_long='1') else '0';
	dataBufferOut(2711) <= dataBufferIn(5185) when (flag_long='1') else '0';
	dataBufferOut(2712) <= dataBufferIn(5928) when (flag_long='1') else '0';
	dataBufferOut(2713) <= dataBufferIn( 527) when (flag_long='1') else '0';
	dataBufferOut(2714) <= dataBufferIn(1270) when (flag_long='1') else '0';
	dataBufferOut(2715) <= dataBufferIn(2013) when (flag_long='1') else '0';
	dataBufferOut(2716) <= dataBufferIn(2756) when (flag_long='1') else '0';
	dataBufferOut(2717) <= dataBufferIn(3499) when (flag_long='1') else '0';
	dataBufferOut(2718) <= dataBufferIn(4242) when (flag_long='1') else '0';
	dataBufferOut(2719) <= dataBufferIn(4985) when (flag_long='1') else '0';
	dataBufferOut(2720) <= dataBufferIn(5728) when (flag_long='1') else '0';
	dataBufferOut(2721) <= dataBufferIn( 327) when (flag_long='1') else '0';
	dataBufferOut(2722) <= dataBufferIn(1070) when (flag_long='1') else '0';
	dataBufferOut(2723) <= dataBufferIn(1813) when (flag_long='1') else '0';
	dataBufferOut(2724) <= dataBufferIn(2556) when (flag_long='1') else '0';
	dataBufferOut(2725) <= dataBufferIn(3299) when (flag_long='1') else '0';
	dataBufferOut(2726) <= dataBufferIn(4042) when (flag_long='1') else '0';
	dataBufferOut(2727) <= dataBufferIn(4785) when (flag_long='1') else '0';
	dataBufferOut(2728) <= dataBufferIn(5528) when (flag_long='1') else '0';
	dataBufferOut(2729) <= dataBufferIn( 127) when (flag_long='1') else '0';
	dataBufferOut(2730) <= dataBufferIn( 870) when (flag_long='1') else '0';
	dataBufferOut(2731) <= dataBufferIn(1613) when (flag_long='1') else '0';
	dataBufferOut(2732) <= dataBufferIn(2356) when (flag_long='1') else '0';
	dataBufferOut(2733) <= dataBufferIn(3099) when (flag_long='1') else '0';
	dataBufferOut(2734) <= dataBufferIn(3842) when (flag_long='1') else '0';
	dataBufferOut(2735) <= dataBufferIn(4585) when (flag_long='1') else '0';
	dataBufferOut(2736) <= dataBufferIn(5328) when (flag_long='1') else '0';
	dataBufferOut(2737) <= dataBufferIn(6071) when (flag_long='1') else '0';
	dataBufferOut(2738) <= dataBufferIn( 670) when (flag_long='1') else '0';
	dataBufferOut(2739) <= dataBufferIn(1413) when (flag_long='1') else '0';
	dataBufferOut(2740) <= dataBufferIn(2156) when (flag_long='1') else '0';
	dataBufferOut(2741) <= dataBufferIn(2899) when (flag_long='1') else '0';
	dataBufferOut(2742) <= dataBufferIn(3642) when (flag_long='1') else '0';
	dataBufferOut(2743) <= dataBufferIn(4385) when (flag_long='1') else '0';
	dataBufferOut(2744) <= dataBufferIn(5128) when (flag_long='1') else '0';
	dataBufferOut(2745) <= dataBufferIn(5871) when (flag_long='1') else '0';
	dataBufferOut(2746) <= dataBufferIn( 470) when (flag_long='1') else '0';
	dataBufferOut(2747) <= dataBufferIn(1213) when (flag_long='1') else '0';
	dataBufferOut(2748) <= dataBufferIn(1956) when (flag_long='1') else '0';
	dataBufferOut(2749) <= dataBufferIn(2699) when (flag_long='1') else '0';
	dataBufferOut(2750) <= dataBufferIn(3442) when (flag_long='1') else '0';
	dataBufferOut(2751) <= dataBufferIn(4185) when (flag_long='1') else '0';
	dataBufferOut(2752) <= dataBufferIn(4928) when (flag_long='1') else '0';
	dataBufferOut(2753) <= dataBufferIn(5671) when (flag_long='1') else '0';
	dataBufferOut(2754) <= dataBufferIn( 270) when (flag_long='1') else '0';
	dataBufferOut(2755) <= dataBufferIn(1013) when (flag_long='1') else '0';
	dataBufferOut(2756) <= dataBufferIn(1756) when (flag_long='1') else '0';
	dataBufferOut(2757) <= dataBufferIn(2499) when (flag_long='1') else '0';
	dataBufferOut(2758) <= dataBufferIn(3242) when (flag_long='1') else '0';
	dataBufferOut(2759) <= dataBufferIn(3985) when (flag_long='1') else '0';
	dataBufferOut(2760) <= dataBufferIn(4728) when (flag_long='1') else '0';
	dataBufferOut(2761) <= dataBufferIn(5471) when (flag_long='1') else '0';
	dataBufferOut(2762) <= dataBufferIn(  70) when (flag_long='1') else '0';
	dataBufferOut(2763) <= dataBufferIn( 813) when (flag_long='1') else '0';
	dataBufferOut(2764) <= dataBufferIn(1556) when (flag_long='1') else '0';
	dataBufferOut(2765) <= dataBufferIn(2299) when (flag_long='1') else '0';
	dataBufferOut(2766) <= dataBufferIn(3042) when (flag_long='1') else '0';
	dataBufferOut(2767) <= dataBufferIn(3785) when (flag_long='1') else '0';
	dataBufferOut(2768) <= dataBufferIn(4528) when (flag_long='1') else '0';
	dataBufferOut(2769) <= dataBufferIn(5271) when (flag_long='1') else '0';
	dataBufferOut(2770) <= dataBufferIn(6014) when (flag_long='1') else '0';
	dataBufferOut(2771) <= dataBufferIn( 613) when (flag_long='1') else '0';
	dataBufferOut(2772) <= dataBufferIn(1356) when (flag_long='1') else '0';
	dataBufferOut(2773) <= dataBufferIn(2099) when (flag_long='1') else '0';
	dataBufferOut(2774) <= dataBufferIn(2842) when (flag_long='1') else '0';
	dataBufferOut(2775) <= dataBufferIn(3585) when (flag_long='1') else '0';
	dataBufferOut(2776) <= dataBufferIn(4328) when (flag_long='1') else '0';
	dataBufferOut(2777) <= dataBufferIn(5071) when (flag_long='1') else '0';
	dataBufferOut(2778) <= dataBufferIn(5814) when (flag_long='1') else '0';
	dataBufferOut(2779) <= dataBufferIn( 413) when (flag_long='1') else '0';
	dataBufferOut(2780) <= dataBufferIn(1156) when (flag_long='1') else '0';
	dataBufferOut(2781) <= dataBufferIn(1899) when (flag_long='1') else '0';
	dataBufferOut(2782) <= dataBufferIn(2642) when (flag_long='1') else '0';
	dataBufferOut(2783) <= dataBufferIn(3385) when (flag_long='1') else '0';
	dataBufferOut(2784) <= dataBufferIn(4128) when (flag_long='1') else '0';
	dataBufferOut(2785) <= dataBufferIn(4871) when (flag_long='1') else '0';
	dataBufferOut(2786) <= dataBufferIn(5614) when (flag_long='1') else '0';
	dataBufferOut(2787) <= dataBufferIn( 213) when (flag_long='1') else '0';
	dataBufferOut(2788) <= dataBufferIn( 956) when (flag_long='1') else '0';
	dataBufferOut(2789) <= dataBufferIn(1699) when (flag_long='1') else '0';
	dataBufferOut(2790) <= dataBufferIn(2442) when (flag_long='1') else '0';
	dataBufferOut(2791) <= dataBufferIn(3185) when (flag_long='1') else '0';
	dataBufferOut(2792) <= dataBufferIn(3928) when (flag_long='1') else '0';
	dataBufferOut(2793) <= dataBufferIn(4671) when (flag_long='1') else '0';
	dataBufferOut(2794) <= dataBufferIn(5414) when (flag_long='1') else '0';
	dataBufferOut(2795) <= dataBufferIn(  13) when (flag_long='1') else '0';
	dataBufferOut(2796) <= dataBufferIn( 756) when (flag_long='1') else '0';
	dataBufferOut(2797) <= dataBufferIn(1499) when (flag_long='1') else '0';
	dataBufferOut(2798) <= dataBufferIn(2242) when (flag_long='1') else '0';
	dataBufferOut(2799) <= dataBufferIn(2985) when (flag_long='1') else '0';
	dataBufferOut(2800) <= dataBufferIn(3728) when (flag_long='1') else '0';
	dataBufferOut(2801) <= dataBufferIn(4471) when (flag_long='1') else '0';
	dataBufferOut(2802) <= dataBufferIn(5214) when (flag_long='1') else '0';
	dataBufferOut(2803) <= dataBufferIn(5957) when (flag_long='1') else '0';
	dataBufferOut(2804) <= dataBufferIn( 556) when (flag_long='1') else '0';
	dataBufferOut(2805) <= dataBufferIn(1299) when (flag_long='1') else '0';
	dataBufferOut(2806) <= dataBufferIn(2042) when (flag_long='1') else '0';
	dataBufferOut(2807) <= dataBufferIn(2785) when (flag_long='1') else '0';
	dataBufferOut(2808) <= dataBufferIn(3528) when (flag_long='1') else '0';
	dataBufferOut(2809) <= dataBufferIn(4271) when (flag_long='1') else '0';
	dataBufferOut(2810) <= dataBufferIn(5014) when (flag_long='1') else '0';
	dataBufferOut(2811) <= dataBufferIn(5757) when (flag_long='1') else '0';
	dataBufferOut(2812) <= dataBufferIn( 356) when (flag_long='1') else '0';
	dataBufferOut(2813) <= dataBufferIn(1099) when (flag_long='1') else '0';
	dataBufferOut(2814) <= dataBufferIn(1842) when (flag_long='1') else '0';
	dataBufferOut(2815) <= dataBufferIn(2585) when (flag_long='1') else '0';
	dataBufferOut(2816) <= dataBufferIn(3328) when (flag_long='1') else '0';
	dataBufferOut(2817) <= dataBufferIn(4071) when (flag_long='1') else '0';
	dataBufferOut(2818) <= dataBufferIn(4814) when (flag_long='1') else '0';
	dataBufferOut(2819) <= dataBufferIn(5557) when (flag_long='1') else '0';
	dataBufferOut(2820) <= dataBufferIn( 156) when (flag_long='1') else '0';
	dataBufferOut(2821) <= dataBufferIn( 899) when (flag_long='1') else '0';
	dataBufferOut(2822) <= dataBufferIn(1642) when (flag_long='1') else '0';
	dataBufferOut(2823) <= dataBufferIn(2385) when (flag_long='1') else '0';
	dataBufferOut(2824) <= dataBufferIn(3128) when (flag_long='1') else '0';
	dataBufferOut(2825) <= dataBufferIn(3871) when (flag_long='1') else '0';
	dataBufferOut(2826) <= dataBufferIn(4614) when (flag_long='1') else '0';
	dataBufferOut(2827) <= dataBufferIn(5357) when (flag_long='1') else '0';
	dataBufferOut(2828) <= dataBufferIn(6100) when (flag_long='1') else '0';
	dataBufferOut(2829) <= dataBufferIn( 699) when (flag_long='1') else '0';
	dataBufferOut(2830) <= dataBufferIn(1442) when (flag_long='1') else '0';
	dataBufferOut(2831) <= dataBufferIn(2185) when (flag_long='1') else '0';
	dataBufferOut(2832) <= dataBufferIn(2928) when (flag_long='1') else '0';
	dataBufferOut(2833) <= dataBufferIn(3671) when (flag_long='1') else '0';
	dataBufferOut(2834) <= dataBufferIn(4414) when (flag_long='1') else '0';
	dataBufferOut(2835) <= dataBufferIn(5157) when (flag_long='1') else '0';
	dataBufferOut(2836) <= dataBufferIn(5900) when (flag_long='1') else '0';
	dataBufferOut(2837) <= dataBufferIn( 499) when (flag_long='1') else '0';
	dataBufferOut(2838) <= dataBufferIn(1242) when (flag_long='1') else '0';
	dataBufferOut(2839) <= dataBufferIn(1985) when (flag_long='1') else '0';
	dataBufferOut(2840) <= dataBufferIn(2728) when (flag_long='1') else '0';
	dataBufferOut(2841) <= dataBufferIn(3471) when (flag_long='1') else '0';
	dataBufferOut(2842) <= dataBufferIn(4214) when (flag_long='1') else '0';
	dataBufferOut(2843) <= dataBufferIn(4957) when (flag_long='1') else '0';
	dataBufferOut(2844) <= dataBufferIn(5700) when (flag_long='1') else '0';
	dataBufferOut(2845) <= dataBufferIn( 299) when (flag_long='1') else '0';
	dataBufferOut(2846) <= dataBufferIn(1042) when (flag_long='1') else '0';
	dataBufferOut(2847) <= dataBufferIn(1785) when (flag_long='1') else '0';
	dataBufferOut(2848) <= dataBufferIn(2528) when (flag_long='1') else '0';
	dataBufferOut(2849) <= dataBufferIn(3271) when (flag_long='1') else '0';
	dataBufferOut(2850) <= dataBufferIn(4014) when (flag_long='1') else '0';
	dataBufferOut(2851) <= dataBufferIn(4757) when (flag_long='1') else '0';
	dataBufferOut(2852) <= dataBufferIn(5500) when (flag_long='1') else '0';
	dataBufferOut(2853) <= dataBufferIn(  99) when (flag_long='1') else '0';
	dataBufferOut(2854) <= dataBufferIn( 842) when (flag_long='1') else '0';
	dataBufferOut(2855) <= dataBufferIn(1585) when (flag_long='1') else '0';
	dataBufferOut(2856) <= dataBufferIn(2328) when (flag_long='1') else '0';
	dataBufferOut(2857) <= dataBufferIn(3071) when (flag_long='1') else '0';
	dataBufferOut(2858) <= dataBufferIn(3814) when (flag_long='1') else '0';
	dataBufferOut(2859) <= dataBufferIn(4557) when (flag_long='1') else '0';
	dataBufferOut(2860) <= dataBufferIn(5300) when (flag_long='1') else '0';
	dataBufferOut(2861) <= dataBufferIn(6043) when (flag_long='1') else '0';
	dataBufferOut(2862) <= dataBufferIn( 642) when (flag_long='1') else '0';
	dataBufferOut(2863) <= dataBufferIn(1385) when (flag_long='1') else '0';
	dataBufferOut(2864) <= dataBufferIn(2128) when (flag_long='1') else '0';
	dataBufferOut(2865) <= dataBufferIn(2871) when (flag_long='1') else '0';
	dataBufferOut(2866) <= dataBufferIn(3614) when (flag_long='1') else '0';
	dataBufferOut(2867) <= dataBufferIn(4357) when (flag_long='1') else '0';
	dataBufferOut(2868) <= dataBufferIn(5100) when (flag_long='1') else '0';
	dataBufferOut(2869) <= dataBufferIn(5843) when (flag_long='1') else '0';
	dataBufferOut(2870) <= dataBufferIn( 442) when (flag_long='1') else '0';
	dataBufferOut(2871) <= dataBufferIn(1185) when (flag_long='1') else '0';
	dataBufferOut(2872) <= dataBufferIn(1928) when (flag_long='1') else '0';
	dataBufferOut(2873) <= dataBufferIn(2671) when (flag_long='1') else '0';
	dataBufferOut(2874) <= dataBufferIn(3414) when (flag_long='1') else '0';
	dataBufferOut(2875) <= dataBufferIn(4157) when (flag_long='1') else '0';
	dataBufferOut(2876) <= dataBufferIn(4900) when (flag_long='1') else '0';
	dataBufferOut(2877) <= dataBufferIn(5643) when (flag_long='1') else '0';
	dataBufferOut(2878) <= dataBufferIn( 242) when (flag_long='1') else '0';
	dataBufferOut(2879) <= dataBufferIn( 985) when (flag_long='1') else '0';
	dataBufferOut(2880) <= dataBufferIn(1728) when (flag_long='1') else '0';
	dataBufferOut(2881) <= dataBufferIn(2471) when (flag_long='1') else '0';
	dataBufferOut(2882) <= dataBufferIn(3214) when (flag_long='1') else '0';
	dataBufferOut(2883) <= dataBufferIn(3957) when (flag_long='1') else '0';
	dataBufferOut(2884) <= dataBufferIn(4700) when (flag_long='1') else '0';
	dataBufferOut(2885) <= dataBufferIn(5443) when (flag_long='1') else '0';
	dataBufferOut(2886) <= dataBufferIn(  42) when (flag_long='1') else '0';
	dataBufferOut(2887) <= dataBufferIn( 785) when (flag_long='1') else '0';
	dataBufferOut(2888) <= dataBufferIn(1528) when (flag_long='1') else '0';
	dataBufferOut(2889) <= dataBufferIn(2271) when (flag_long='1') else '0';
	dataBufferOut(2890) <= dataBufferIn(3014) when (flag_long='1') else '0';
	dataBufferOut(2891) <= dataBufferIn(3757) when (flag_long='1') else '0';
	dataBufferOut(2892) <= dataBufferIn(4500) when (flag_long='1') else '0';
	dataBufferOut(2893) <= dataBufferIn(5243) when (flag_long='1') else '0';
	dataBufferOut(2894) <= dataBufferIn(5986) when (flag_long='1') else '0';
	dataBufferOut(2895) <= dataBufferIn( 585) when (flag_long='1') else '0';
	dataBufferOut(2896) <= dataBufferIn(1328) when (flag_long='1') else '0';
	dataBufferOut(2897) <= dataBufferIn(2071) when (flag_long='1') else '0';
	dataBufferOut(2898) <= dataBufferIn(2814) when (flag_long='1') else '0';
	dataBufferOut(2899) <= dataBufferIn(3557) when (flag_long='1') else '0';
	dataBufferOut(2900) <= dataBufferIn(4300) when (flag_long='1') else '0';
	dataBufferOut(2901) <= dataBufferIn(5043) when (flag_long='1') else '0';
	dataBufferOut(2902) <= dataBufferIn(5786) when (flag_long='1') else '0';
	dataBufferOut(2903) <= dataBufferIn( 385) when (flag_long='1') else '0';
	dataBufferOut(2904) <= dataBufferIn(1128) when (flag_long='1') else '0';
	dataBufferOut(2905) <= dataBufferIn(1871) when (flag_long='1') else '0';
	dataBufferOut(2906) <= dataBufferIn(2614) when (flag_long='1') else '0';
	dataBufferOut(2907) <= dataBufferIn(3357) when (flag_long='1') else '0';
	dataBufferOut(2908) <= dataBufferIn(4100) when (flag_long='1') else '0';
	dataBufferOut(2909) <= dataBufferIn(4843) when (flag_long='1') else '0';
	dataBufferOut(2910) <= dataBufferIn(5586) when (flag_long='1') else '0';
	dataBufferOut(2911) <= dataBufferIn( 185) when (flag_long='1') else '0';
	dataBufferOut(2912) <= dataBufferIn( 928) when (flag_long='1') else '0';
	dataBufferOut(2913) <= dataBufferIn(1671) when (flag_long='1') else '0';
	dataBufferOut(2914) <= dataBufferIn(2414) when (flag_long='1') else '0';
	dataBufferOut(2915) <= dataBufferIn(3157) when (flag_long='1') else '0';
	dataBufferOut(2916) <= dataBufferIn(3900) when (flag_long='1') else '0';
	dataBufferOut(2917) <= dataBufferIn(4643) when (flag_long='1') else '0';
	dataBufferOut(2918) <= dataBufferIn(5386) when (flag_long='1') else '0';
	dataBufferOut(2919) <= dataBufferIn(6129) when (flag_long='1') else '0';
	dataBufferOut(2920) <= dataBufferIn( 728) when (flag_long='1') else '0';
	dataBufferOut(2921) <= dataBufferIn(1471) when (flag_long='1') else '0';
	dataBufferOut(2922) <= dataBufferIn(2214) when (flag_long='1') else '0';
	dataBufferOut(2923) <= dataBufferIn(2957) when (flag_long='1') else '0';
	dataBufferOut(2924) <= dataBufferIn(3700) when (flag_long='1') else '0';
	dataBufferOut(2925) <= dataBufferIn(4443) when (flag_long='1') else '0';
	dataBufferOut(2926) <= dataBufferIn(5186) when (flag_long='1') else '0';
	dataBufferOut(2927) <= dataBufferIn(5929) when (flag_long='1') else '0';
	dataBufferOut(2928) <= dataBufferIn( 528) when (flag_long='1') else '0';
	dataBufferOut(2929) <= dataBufferIn(1271) when (flag_long='1') else '0';
	dataBufferOut(2930) <= dataBufferIn(2014) when (flag_long='1') else '0';
	dataBufferOut(2931) <= dataBufferIn(2757) when (flag_long='1') else '0';
	dataBufferOut(2932) <= dataBufferIn(3500) when (flag_long='1') else '0';
	dataBufferOut(2933) <= dataBufferIn(4243) when (flag_long='1') else '0';
	dataBufferOut(2934) <= dataBufferIn(4986) when (flag_long='1') else '0';
	dataBufferOut(2935) <= dataBufferIn(5729) when (flag_long='1') else '0';
	dataBufferOut(2936) <= dataBufferIn( 328) when (flag_long='1') else '0';
	dataBufferOut(2937) <= dataBufferIn(1071) when (flag_long='1') else '0';
	dataBufferOut(2938) <= dataBufferIn(1814) when (flag_long='1') else '0';
	dataBufferOut(2939) <= dataBufferIn(2557) when (flag_long='1') else '0';
	dataBufferOut(2940) <= dataBufferIn(3300) when (flag_long='1') else '0';
	dataBufferOut(2941) <= dataBufferIn(4043) when (flag_long='1') else '0';
	dataBufferOut(2942) <= dataBufferIn(4786) when (flag_long='1') else '0';
	dataBufferOut(2943) <= dataBufferIn(5529) when (flag_long='1') else '0';
	dataBufferOut(2944) <= dataBufferIn( 128) when (flag_long='1') else '0';
	dataBufferOut(2945) <= dataBufferIn( 871) when (flag_long='1') else '0';
	dataBufferOut(2946) <= dataBufferIn(1614) when (flag_long='1') else '0';
	dataBufferOut(2947) <= dataBufferIn(2357) when (flag_long='1') else '0';
	dataBufferOut(2948) <= dataBufferIn(3100) when (flag_long='1') else '0';
	dataBufferOut(2949) <= dataBufferIn(3843) when (flag_long='1') else '0';
	dataBufferOut(2950) <= dataBufferIn(4586) when (flag_long='1') else '0';
	dataBufferOut(2951) <= dataBufferIn(5329) when (flag_long='1') else '0';
	dataBufferOut(2952) <= dataBufferIn(6072) when (flag_long='1') else '0';
	dataBufferOut(2953) <= dataBufferIn( 671) when (flag_long='1') else '0';
	dataBufferOut(2954) <= dataBufferIn(1414) when (flag_long='1') else '0';
	dataBufferOut(2955) <= dataBufferIn(2157) when (flag_long='1') else '0';
	dataBufferOut(2956) <= dataBufferIn(2900) when (flag_long='1') else '0';
	dataBufferOut(2957) <= dataBufferIn(3643) when (flag_long='1') else '0';
	dataBufferOut(2958) <= dataBufferIn(4386) when (flag_long='1') else '0';
	dataBufferOut(2959) <= dataBufferIn(5129) when (flag_long='1') else '0';
	dataBufferOut(2960) <= dataBufferIn(5872) when (flag_long='1') else '0';
	dataBufferOut(2961) <= dataBufferIn( 471) when (flag_long='1') else '0';
	dataBufferOut(2962) <= dataBufferIn(1214) when (flag_long='1') else '0';
	dataBufferOut(2963) <= dataBufferIn(1957) when (flag_long='1') else '0';
	dataBufferOut(2964) <= dataBufferIn(2700) when (flag_long='1') else '0';
	dataBufferOut(2965) <= dataBufferIn(3443) when (flag_long='1') else '0';
	dataBufferOut(2966) <= dataBufferIn(4186) when (flag_long='1') else '0';
	dataBufferOut(2967) <= dataBufferIn(4929) when (flag_long='1') else '0';
	dataBufferOut(2968) <= dataBufferIn(5672) when (flag_long='1') else '0';
	dataBufferOut(2969) <= dataBufferIn( 271) when (flag_long='1') else '0';
	dataBufferOut(2970) <= dataBufferIn(1014) when (flag_long='1') else '0';
	dataBufferOut(2971) <= dataBufferIn(1757) when (flag_long='1') else '0';
	dataBufferOut(2972) <= dataBufferIn(2500) when (flag_long='1') else '0';
	dataBufferOut(2973) <= dataBufferIn(3243) when (flag_long='1') else '0';
	dataBufferOut(2974) <= dataBufferIn(3986) when (flag_long='1') else '0';
	dataBufferOut(2975) <= dataBufferIn(4729) when (flag_long='1') else '0';
	dataBufferOut(2976) <= dataBufferIn(5472) when (flag_long='1') else '0';
	dataBufferOut(2977) <= dataBufferIn(  71) when (flag_long='1') else '0';
	dataBufferOut(2978) <= dataBufferIn( 814) when (flag_long='1') else '0';
	dataBufferOut(2979) <= dataBufferIn(1557) when (flag_long='1') else '0';
	dataBufferOut(2980) <= dataBufferIn(2300) when (flag_long='1') else '0';
	dataBufferOut(2981) <= dataBufferIn(3043) when (flag_long='1') else '0';
	dataBufferOut(2982) <= dataBufferIn(3786) when (flag_long='1') else '0';
	dataBufferOut(2983) <= dataBufferIn(4529) when (flag_long='1') else '0';
	dataBufferOut(2984) <= dataBufferIn(5272) when (flag_long='1') else '0';
	dataBufferOut(2985) <= dataBufferIn(6015) when (flag_long='1') else '0';
	dataBufferOut(2986) <= dataBufferIn( 614) when (flag_long='1') else '0';
	dataBufferOut(2987) <= dataBufferIn(1357) when (flag_long='1') else '0';
	dataBufferOut(2988) <= dataBufferIn(2100) when (flag_long='1') else '0';
	dataBufferOut(2989) <= dataBufferIn(2843) when (flag_long='1') else '0';
	dataBufferOut(2990) <= dataBufferIn(3586) when (flag_long='1') else '0';
	dataBufferOut(2991) <= dataBufferIn(4329) when (flag_long='1') else '0';
	dataBufferOut(2992) <= dataBufferIn(5072) when (flag_long='1') else '0';
	dataBufferOut(2993) <= dataBufferIn(5815) when (flag_long='1') else '0';
	dataBufferOut(2994) <= dataBufferIn( 414) when (flag_long='1') else '0';
	dataBufferOut(2995) <= dataBufferIn(1157) when (flag_long='1') else '0';
	dataBufferOut(2996) <= dataBufferIn(1900) when (flag_long='1') else '0';
	dataBufferOut(2997) <= dataBufferIn(2643) when (flag_long='1') else '0';
	dataBufferOut(2998) <= dataBufferIn(3386) when (flag_long='1') else '0';
	dataBufferOut(2999) <= dataBufferIn(4129) when (flag_long='1') else '0';
	dataBufferOut(3000) <= dataBufferIn(4872) when (flag_long='1') else '0';
	dataBufferOut(3001) <= dataBufferIn(5615) when (flag_long='1') else '0';
	dataBufferOut(3002) <= dataBufferIn( 214) when (flag_long='1') else '0';
	dataBufferOut(3003) <= dataBufferIn( 957) when (flag_long='1') else '0';
	dataBufferOut(3004) <= dataBufferIn(1700) when (flag_long='1') else '0';
	dataBufferOut(3005) <= dataBufferIn(2443) when (flag_long='1') else '0';
	dataBufferOut(3006) <= dataBufferIn(3186) when (flag_long='1') else '0';
	dataBufferOut(3007) <= dataBufferIn(3929) when (flag_long='1') else '0';
	dataBufferOut(3008) <= dataBufferIn(4672) when (flag_long='1') else '0';
	dataBufferOut(3009) <= dataBufferIn(5415) when (flag_long='1') else '0';
	dataBufferOut(3010) <= dataBufferIn(  14) when (flag_long='1') else '0';
	dataBufferOut(3011) <= dataBufferIn( 757) when (flag_long='1') else '0';
	dataBufferOut(3012) <= dataBufferIn(1500) when (flag_long='1') else '0';
	dataBufferOut(3013) <= dataBufferIn(2243) when (flag_long='1') else '0';
	dataBufferOut(3014) <= dataBufferIn(2986) when (flag_long='1') else '0';
	dataBufferOut(3015) <= dataBufferIn(3729) when (flag_long='1') else '0';
	dataBufferOut(3016) <= dataBufferIn(4472) when (flag_long='1') else '0';
	dataBufferOut(3017) <= dataBufferIn(5215) when (flag_long='1') else '0';
	dataBufferOut(3018) <= dataBufferIn(5958) when (flag_long='1') else '0';
	dataBufferOut(3019) <= dataBufferIn( 557) when (flag_long='1') else '0';
	dataBufferOut(3020) <= dataBufferIn(1300) when (flag_long='1') else '0';
	dataBufferOut(3021) <= dataBufferIn(2043) when (flag_long='1') else '0';
	dataBufferOut(3022) <= dataBufferIn(2786) when (flag_long='1') else '0';
	dataBufferOut(3023) <= dataBufferIn(3529) when (flag_long='1') else '0';
	dataBufferOut(3024) <= dataBufferIn(4272) when (flag_long='1') else '0';
	dataBufferOut(3025) <= dataBufferIn(5015) when (flag_long='1') else '0';
	dataBufferOut(3026) <= dataBufferIn(5758) when (flag_long='1') else '0';
	dataBufferOut(3027) <= dataBufferIn( 357) when (flag_long='1') else '0';
	dataBufferOut(3028) <= dataBufferIn(1100) when (flag_long='1') else '0';
	dataBufferOut(3029) <= dataBufferIn(1843) when (flag_long='1') else '0';
	dataBufferOut(3030) <= dataBufferIn(2586) when (flag_long='1') else '0';
	dataBufferOut(3031) <= dataBufferIn(3329) when (flag_long='1') else '0';
	dataBufferOut(3032) <= dataBufferIn(4072) when (flag_long='1') else '0';
	dataBufferOut(3033) <= dataBufferIn(4815) when (flag_long='1') else '0';
	dataBufferOut(3034) <= dataBufferIn(5558) when (flag_long='1') else '0';
	dataBufferOut(3035) <= dataBufferIn( 157) when (flag_long='1') else '0';
	dataBufferOut(3036) <= dataBufferIn( 900) when (flag_long='1') else '0';
	dataBufferOut(3037) <= dataBufferIn(1643) when (flag_long='1') else '0';
	dataBufferOut(3038) <= dataBufferIn(2386) when (flag_long='1') else '0';
	dataBufferOut(3039) <= dataBufferIn(3129) when (flag_long='1') else '0';
	dataBufferOut(3040) <= dataBufferIn(3872) when (flag_long='1') else '0';
	dataBufferOut(3041) <= dataBufferIn(4615) when (flag_long='1') else '0';
	dataBufferOut(3042) <= dataBufferIn(5358) when (flag_long='1') else '0';
	dataBufferOut(3043) <= dataBufferIn(6101) when (flag_long='1') else '0';
	dataBufferOut(3044) <= dataBufferIn( 700) when (flag_long='1') else '0';
	dataBufferOut(3045) <= dataBufferIn(1443) when (flag_long='1') else '0';
	dataBufferOut(3046) <= dataBufferIn(2186) when (flag_long='1') else '0';
	dataBufferOut(3047) <= dataBufferIn(2929) when (flag_long='1') else '0';
	dataBufferOut(3048) <= dataBufferIn(3672) when (flag_long='1') else '0';
	dataBufferOut(3049) <= dataBufferIn(4415) when (flag_long='1') else '0';
	dataBufferOut(3050) <= dataBufferIn(5158) when (flag_long='1') else '0';
	dataBufferOut(3051) <= dataBufferIn(5901) when (flag_long='1') else '0';
	dataBufferOut(3052) <= dataBufferIn( 500) when (flag_long='1') else '0';
	dataBufferOut(3053) <= dataBufferIn(1243) when (flag_long='1') else '0';
	dataBufferOut(3054) <= dataBufferIn(1986) when (flag_long='1') else '0';
	dataBufferOut(3055) <= dataBufferIn(2729) when (flag_long='1') else '0';
	dataBufferOut(3056) <= dataBufferIn(3472) when (flag_long='1') else '0';
	dataBufferOut(3057) <= dataBufferIn(4215) when (flag_long='1') else '0';
	dataBufferOut(3058) <= dataBufferIn(4958) when (flag_long='1') else '0';
	dataBufferOut(3059) <= dataBufferIn(5701) when (flag_long='1') else '0';
	dataBufferOut(3060) <= dataBufferIn( 300) when (flag_long='1') else '0';
	dataBufferOut(3061) <= dataBufferIn(1043) when (flag_long='1') else '0';
	dataBufferOut(3062) <= dataBufferIn(1786) when (flag_long='1') else '0';
	dataBufferOut(3063) <= dataBufferIn(2529) when (flag_long='1') else '0';
	dataBufferOut(3064) <= dataBufferIn(3272) when (flag_long='1') else '0';
	dataBufferOut(3065) <= dataBufferIn(4015) when (flag_long='1') else '0';
	dataBufferOut(3066) <= dataBufferIn(4758) when (flag_long='1') else '0';
	dataBufferOut(3067) <= dataBufferIn(5501) when (flag_long='1') else '0';
	dataBufferOut(3068) <= dataBufferIn( 100) when (flag_long='1') else '0';
	dataBufferOut(3069) <= dataBufferIn( 843) when (flag_long='1') else '0';
	dataBufferOut(3070) <= dataBufferIn(1586) when (flag_long='1') else '0';
	dataBufferOut(3071) <= dataBufferIn(2329) when (flag_long='1') else '0';
	dataBufferOut(3072) <= dataBufferIn(3072) when (flag_long='1') else '0';
	dataBufferOut(3073) <= dataBufferIn(3815) when (flag_long='1') else '0';
	dataBufferOut(3074) <= dataBufferIn(4558) when (flag_long='1') else '0';
	dataBufferOut(3075) <= dataBufferIn(5301) when (flag_long='1') else '0';
	dataBufferOut(3076) <= dataBufferIn(6044) when (flag_long='1') else '0';
	dataBufferOut(3077) <= dataBufferIn( 643) when (flag_long='1') else '0';
	dataBufferOut(3078) <= dataBufferIn(1386) when (flag_long='1') else '0';
	dataBufferOut(3079) <= dataBufferIn(2129) when (flag_long='1') else '0';
	dataBufferOut(3080) <= dataBufferIn(2872) when (flag_long='1') else '0';
	dataBufferOut(3081) <= dataBufferIn(3615) when (flag_long='1') else '0';
	dataBufferOut(3082) <= dataBufferIn(4358) when (flag_long='1') else '0';
	dataBufferOut(3083) <= dataBufferIn(5101) when (flag_long='1') else '0';
	dataBufferOut(3084) <= dataBufferIn(5844) when (flag_long='1') else '0';
	dataBufferOut(3085) <= dataBufferIn( 443) when (flag_long='1') else '0';
	dataBufferOut(3086) <= dataBufferIn(1186) when (flag_long='1') else '0';
	dataBufferOut(3087) <= dataBufferIn(1929) when (flag_long='1') else '0';
	dataBufferOut(3088) <= dataBufferIn(2672) when (flag_long='1') else '0';
	dataBufferOut(3089) <= dataBufferIn(3415) when (flag_long='1') else '0';
	dataBufferOut(3090) <= dataBufferIn(4158) when (flag_long='1') else '0';
	dataBufferOut(3091) <= dataBufferIn(4901) when (flag_long='1') else '0';
	dataBufferOut(3092) <= dataBufferIn(5644) when (flag_long='1') else '0';
	dataBufferOut(3093) <= dataBufferIn( 243) when (flag_long='1') else '0';
	dataBufferOut(3094) <= dataBufferIn( 986) when (flag_long='1') else '0';
	dataBufferOut(3095) <= dataBufferIn(1729) when (flag_long='1') else '0';
	dataBufferOut(3096) <= dataBufferIn(2472) when (flag_long='1') else '0';
	dataBufferOut(3097) <= dataBufferIn(3215) when (flag_long='1') else '0';
	dataBufferOut(3098) <= dataBufferIn(3958) when (flag_long='1') else '0';
	dataBufferOut(3099) <= dataBufferIn(4701) when (flag_long='1') else '0';
	dataBufferOut(3100) <= dataBufferIn(5444) when (flag_long='1') else '0';
	dataBufferOut(3101) <= dataBufferIn(  43) when (flag_long='1') else '0';
	dataBufferOut(3102) <= dataBufferIn( 786) when (flag_long='1') else '0';
	dataBufferOut(3103) <= dataBufferIn(1529) when (flag_long='1') else '0';
	dataBufferOut(3104) <= dataBufferIn(2272) when (flag_long='1') else '0';
	dataBufferOut(3105) <= dataBufferIn(3015) when (flag_long='1') else '0';
	dataBufferOut(3106) <= dataBufferIn(3758) when (flag_long='1') else '0';
	dataBufferOut(3107) <= dataBufferIn(4501) when (flag_long='1') else '0';
	dataBufferOut(3108) <= dataBufferIn(5244) when (flag_long='1') else '0';
	dataBufferOut(3109) <= dataBufferIn(5987) when (flag_long='1') else '0';
	dataBufferOut(3110) <= dataBufferIn( 586) when (flag_long='1') else '0';
	dataBufferOut(3111) <= dataBufferIn(1329) when (flag_long='1') else '0';
	dataBufferOut(3112) <= dataBufferIn(2072) when (flag_long='1') else '0';
	dataBufferOut(3113) <= dataBufferIn(2815) when (flag_long='1') else '0';
	dataBufferOut(3114) <= dataBufferIn(3558) when (flag_long='1') else '0';
	dataBufferOut(3115) <= dataBufferIn(4301) when (flag_long='1') else '0';
	dataBufferOut(3116) <= dataBufferIn(5044) when (flag_long='1') else '0';
	dataBufferOut(3117) <= dataBufferIn(5787) when (flag_long='1') else '0';
	dataBufferOut(3118) <= dataBufferIn( 386) when (flag_long='1') else '0';
	dataBufferOut(3119) <= dataBufferIn(1129) when (flag_long='1') else '0';
	dataBufferOut(3120) <= dataBufferIn(1872) when (flag_long='1') else '0';
	dataBufferOut(3121) <= dataBufferIn(2615) when (flag_long='1') else '0';
	dataBufferOut(3122) <= dataBufferIn(3358) when (flag_long='1') else '0';
	dataBufferOut(3123) <= dataBufferIn(4101) when (flag_long='1') else '0';
	dataBufferOut(3124) <= dataBufferIn(4844) when (flag_long='1') else '0';
	dataBufferOut(3125) <= dataBufferIn(5587) when (flag_long='1') else '0';
	dataBufferOut(3126) <= dataBufferIn( 186) when (flag_long='1') else '0';
	dataBufferOut(3127) <= dataBufferIn( 929) when (flag_long='1') else '0';
	dataBufferOut(3128) <= dataBufferIn(1672) when (flag_long='1') else '0';
	dataBufferOut(3129) <= dataBufferIn(2415) when (flag_long='1') else '0';
	dataBufferOut(3130) <= dataBufferIn(3158) when (flag_long='1') else '0';
	dataBufferOut(3131) <= dataBufferIn(3901) when (flag_long='1') else '0';
	dataBufferOut(3132) <= dataBufferIn(4644) when (flag_long='1') else '0';
	dataBufferOut(3133) <= dataBufferIn(5387) when (flag_long='1') else '0';
	dataBufferOut(3134) <= dataBufferIn(6130) when (flag_long='1') else '0';
	dataBufferOut(3135) <= dataBufferIn( 729) when (flag_long='1') else '0';
	dataBufferOut(3136) <= dataBufferIn(1472) when (flag_long='1') else '0';
	dataBufferOut(3137) <= dataBufferIn(2215) when (flag_long='1') else '0';
	dataBufferOut(3138) <= dataBufferIn(2958) when (flag_long='1') else '0';
	dataBufferOut(3139) <= dataBufferIn(3701) when (flag_long='1') else '0';
	dataBufferOut(3140) <= dataBufferIn(4444) when (flag_long='1') else '0';
	dataBufferOut(3141) <= dataBufferIn(5187) when (flag_long='1') else '0';
	dataBufferOut(3142) <= dataBufferIn(5930) when (flag_long='1') else '0';
	dataBufferOut(3143) <= dataBufferIn( 529) when (flag_long='1') else '0';
	dataBufferOut(3144) <= dataBufferIn(1272) when (flag_long='1') else '0';
	dataBufferOut(3145) <= dataBufferIn(2015) when (flag_long='1') else '0';
	dataBufferOut(3146) <= dataBufferIn(2758) when (flag_long='1') else '0';
	dataBufferOut(3147) <= dataBufferIn(3501) when (flag_long='1') else '0';
	dataBufferOut(3148) <= dataBufferIn(4244) when (flag_long='1') else '0';
	dataBufferOut(3149) <= dataBufferIn(4987) when (flag_long='1') else '0';
	dataBufferOut(3150) <= dataBufferIn(5730) when (flag_long='1') else '0';
	dataBufferOut(3151) <= dataBufferIn( 329) when (flag_long='1') else '0';
	dataBufferOut(3152) <= dataBufferIn(1072) when (flag_long='1') else '0';
	dataBufferOut(3153) <= dataBufferIn(1815) when (flag_long='1') else '0';
	dataBufferOut(3154) <= dataBufferIn(2558) when (flag_long='1') else '0';
	dataBufferOut(3155) <= dataBufferIn(3301) when (flag_long='1') else '0';
	dataBufferOut(3156) <= dataBufferIn(4044) when (flag_long='1') else '0';
	dataBufferOut(3157) <= dataBufferIn(4787) when (flag_long='1') else '0';
	dataBufferOut(3158) <= dataBufferIn(5530) when (flag_long='1') else '0';
	dataBufferOut(3159) <= dataBufferIn( 129) when (flag_long='1') else '0';
	dataBufferOut(3160) <= dataBufferIn( 872) when (flag_long='1') else '0';
	dataBufferOut(3161) <= dataBufferIn(1615) when (flag_long='1') else '0';
	dataBufferOut(3162) <= dataBufferIn(2358) when (flag_long='1') else '0';
	dataBufferOut(3163) <= dataBufferIn(3101) when (flag_long='1') else '0';
	dataBufferOut(3164) <= dataBufferIn(3844) when (flag_long='1') else '0';
	dataBufferOut(3165) <= dataBufferIn(4587) when (flag_long='1') else '0';
	dataBufferOut(3166) <= dataBufferIn(5330) when (flag_long='1') else '0';
	dataBufferOut(3167) <= dataBufferIn(6073) when (flag_long='1') else '0';
	dataBufferOut(3168) <= dataBufferIn( 672) when (flag_long='1') else '0';
	dataBufferOut(3169) <= dataBufferIn(1415) when (flag_long='1') else '0';
	dataBufferOut(3170) <= dataBufferIn(2158) when (flag_long='1') else '0';
	dataBufferOut(3171) <= dataBufferIn(2901) when (flag_long='1') else '0';
	dataBufferOut(3172) <= dataBufferIn(3644) when (flag_long='1') else '0';
	dataBufferOut(3173) <= dataBufferIn(4387) when (flag_long='1') else '0';
	dataBufferOut(3174) <= dataBufferIn(5130) when (flag_long='1') else '0';
	dataBufferOut(3175) <= dataBufferIn(5873) when (flag_long='1') else '0';
	dataBufferOut(3176) <= dataBufferIn( 472) when (flag_long='1') else '0';
	dataBufferOut(3177) <= dataBufferIn(1215) when (flag_long='1') else '0';
	dataBufferOut(3178) <= dataBufferIn(1958) when (flag_long='1') else '0';
	dataBufferOut(3179) <= dataBufferIn(2701) when (flag_long='1') else '0';
	dataBufferOut(3180) <= dataBufferIn(3444) when (flag_long='1') else '0';
	dataBufferOut(3181) <= dataBufferIn(4187) when (flag_long='1') else '0';
	dataBufferOut(3182) <= dataBufferIn(4930) when (flag_long='1') else '0';
	dataBufferOut(3183) <= dataBufferIn(5673) when (flag_long='1') else '0';
	dataBufferOut(3184) <= dataBufferIn( 272) when (flag_long='1') else '0';
	dataBufferOut(3185) <= dataBufferIn(1015) when (flag_long='1') else '0';
	dataBufferOut(3186) <= dataBufferIn(1758) when (flag_long='1') else '0';
	dataBufferOut(3187) <= dataBufferIn(2501) when (flag_long='1') else '0';
	dataBufferOut(3188) <= dataBufferIn(3244) when (flag_long='1') else '0';
	dataBufferOut(3189) <= dataBufferIn(3987) when (flag_long='1') else '0';
	dataBufferOut(3190) <= dataBufferIn(4730) when (flag_long='1') else '0';
	dataBufferOut(3191) <= dataBufferIn(5473) when (flag_long='1') else '0';
	dataBufferOut(3192) <= dataBufferIn(  72) when (flag_long='1') else '0';
	dataBufferOut(3193) <= dataBufferIn( 815) when (flag_long='1') else '0';
	dataBufferOut(3194) <= dataBufferIn(1558) when (flag_long='1') else '0';
	dataBufferOut(3195) <= dataBufferIn(2301) when (flag_long='1') else '0';
	dataBufferOut(3196) <= dataBufferIn(3044) when (flag_long='1') else '0';
	dataBufferOut(3197) <= dataBufferIn(3787) when (flag_long='1') else '0';
	dataBufferOut(3198) <= dataBufferIn(4530) when (flag_long='1') else '0';
	dataBufferOut(3199) <= dataBufferIn(5273) when (flag_long='1') else '0';
	dataBufferOut(3200) <= dataBufferIn(6016) when (flag_long='1') else '0';
	dataBufferOut(3201) <= dataBufferIn( 615) when (flag_long='1') else '0';
	dataBufferOut(3202) <= dataBufferIn(1358) when (flag_long='1') else '0';
	dataBufferOut(3203) <= dataBufferIn(2101) when (flag_long='1') else '0';
	dataBufferOut(3204) <= dataBufferIn(2844) when (flag_long='1') else '0';
	dataBufferOut(3205) <= dataBufferIn(3587) when (flag_long='1') else '0';
	dataBufferOut(3206) <= dataBufferIn(4330) when (flag_long='1') else '0';
	dataBufferOut(3207) <= dataBufferIn(5073) when (flag_long='1') else '0';
	dataBufferOut(3208) <= dataBufferIn(5816) when (flag_long='1') else '0';
	dataBufferOut(3209) <= dataBufferIn( 415) when (flag_long='1') else '0';
	dataBufferOut(3210) <= dataBufferIn(1158) when (flag_long='1') else '0';
	dataBufferOut(3211) <= dataBufferIn(1901) when (flag_long='1') else '0';
	dataBufferOut(3212) <= dataBufferIn(2644) when (flag_long='1') else '0';
	dataBufferOut(3213) <= dataBufferIn(3387) when (flag_long='1') else '0';
	dataBufferOut(3214) <= dataBufferIn(4130) when (flag_long='1') else '0';
	dataBufferOut(3215) <= dataBufferIn(4873) when (flag_long='1') else '0';
	dataBufferOut(3216) <= dataBufferIn(5616) when (flag_long='1') else '0';
	dataBufferOut(3217) <= dataBufferIn( 215) when (flag_long='1') else '0';
	dataBufferOut(3218) <= dataBufferIn( 958) when (flag_long='1') else '0';
	dataBufferOut(3219) <= dataBufferIn(1701) when (flag_long='1') else '0';
	dataBufferOut(3220) <= dataBufferIn(2444) when (flag_long='1') else '0';
	dataBufferOut(3221) <= dataBufferIn(3187) when (flag_long='1') else '0';
	dataBufferOut(3222) <= dataBufferIn(3930) when (flag_long='1') else '0';
	dataBufferOut(3223) <= dataBufferIn(4673) when (flag_long='1') else '0';
	dataBufferOut(3224) <= dataBufferIn(5416) when (flag_long='1') else '0';
	dataBufferOut(3225) <= dataBufferIn(  15) when (flag_long='1') else '0';
	dataBufferOut(3226) <= dataBufferIn( 758) when (flag_long='1') else '0';
	dataBufferOut(3227) <= dataBufferIn(1501) when (flag_long='1') else '0';
	dataBufferOut(3228) <= dataBufferIn(2244) when (flag_long='1') else '0';
	dataBufferOut(3229) <= dataBufferIn(2987) when (flag_long='1') else '0';
	dataBufferOut(3230) <= dataBufferIn(3730) when (flag_long='1') else '0';
	dataBufferOut(3231) <= dataBufferIn(4473) when (flag_long='1') else '0';
	dataBufferOut(3232) <= dataBufferIn(5216) when (flag_long='1') else '0';
	dataBufferOut(3233) <= dataBufferIn(5959) when (flag_long='1') else '0';
	dataBufferOut(3234) <= dataBufferIn( 558) when (flag_long='1') else '0';
	dataBufferOut(3235) <= dataBufferIn(1301) when (flag_long='1') else '0';
	dataBufferOut(3236) <= dataBufferIn(2044) when (flag_long='1') else '0';
	dataBufferOut(3237) <= dataBufferIn(2787) when (flag_long='1') else '0';
	dataBufferOut(3238) <= dataBufferIn(3530) when (flag_long='1') else '0';
	dataBufferOut(3239) <= dataBufferIn(4273) when (flag_long='1') else '0';
	dataBufferOut(3240) <= dataBufferIn(5016) when (flag_long='1') else '0';
	dataBufferOut(3241) <= dataBufferIn(5759) when (flag_long='1') else '0';
	dataBufferOut(3242) <= dataBufferIn( 358) when (flag_long='1') else '0';
	dataBufferOut(3243) <= dataBufferIn(1101) when (flag_long='1') else '0';
	dataBufferOut(3244) <= dataBufferIn(1844) when (flag_long='1') else '0';
	dataBufferOut(3245) <= dataBufferIn(2587) when (flag_long='1') else '0';
	dataBufferOut(3246) <= dataBufferIn(3330) when (flag_long='1') else '0';
	dataBufferOut(3247) <= dataBufferIn(4073) when (flag_long='1') else '0';
	dataBufferOut(3248) <= dataBufferIn(4816) when (flag_long='1') else '0';
	dataBufferOut(3249) <= dataBufferIn(5559) when (flag_long='1') else '0';
	dataBufferOut(3250) <= dataBufferIn( 158) when (flag_long='1') else '0';
	dataBufferOut(3251) <= dataBufferIn( 901) when (flag_long='1') else '0';
	dataBufferOut(3252) <= dataBufferIn(1644) when (flag_long='1') else '0';
	dataBufferOut(3253) <= dataBufferIn(2387) when (flag_long='1') else '0';
	dataBufferOut(3254) <= dataBufferIn(3130) when (flag_long='1') else '0';
	dataBufferOut(3255) <= dataBufferIn(3873) when (flag_long='1') else '0';
	dataBufferOut(3256) <= dataBufferIn(4616) when (flag_long='1') else '0';
	dataBufferOut(3257) <= dataBufferIn(5359) when (flag_long='1') else '0';
	dataBufferOut(3258) <= dataBufferIn(6102) when (flag_long='1') else '0';
	dataBufferOut(3259) <= dataBufferIn( 701) when (flag_long='1') else '0';
	dataBufferOut(3260) <= dataBufferIn(1444) when (flag_long='1') else '0';
	dataBufferOut(3261) <= dataBufferIn(2187) when (flag_long='1') else '0';
	dataBufferOut(3262) <= dataBufferIn(2930) when (flag_long='1') else '0';
	dataBufferOut(3263) <= dataBufferIn(3673) when (flag_long='1') else '0';
	dataBufferOut(3264) <= dataBufferIn(4416) when (flag_long='1') else '0';
	dataBufferOut(3265) <= dataBufferIn(5159) when (flag_long='1') else '0';
	dataBufferOut(3266) <= dataBufferIn(5902) when (flag_long='1') else '0';
	dataBufferOut(3267) <= dataBufferIn( 501) when (flag_long='1') else '0';
	dataBufferOut(3268) <= dataBufferIn(1244) when (flag_long='1') else '0';
	dataBufferOut(3269) <= dataBufferIn(1987) when (flag_long='1') else '0';
	dataBufferOut(3270) <= dataBufferIn(2730) when (flag_long='1') else '0';
	dataBufferOut(3271) <= dataBufferIn(3473) when (flag_long='1') else '0';
	dataBufferOut(3272) <= dataBufferIn(4216) when (flag_long='1') else '0';
	dataBufferOut(3273) <= dataBufferIn(4959) when (flag_long='1') else '0';
	dataBufferOut(3274) <= dataBufferIn(5702) when (flag_long='1') else '0';
	dataBufferOut(3275) <= dataBufferIn( 301) when (flag_long='1') else '0';
	dataBufferOut(3276) <= dataBufferIn(1044) when (flag_long='1') else '0';
	dataBufferOut(3277) <= dataBufferIn(1787) when (flag_long='1') else '0';
	dataBufferOut(3278) <= dataBufferIn(2530) when (flag_long='1') else '0';
	dataBufferOut(3279) <= dataBufferIn(3273) when (flag_long='1') else '0';
	dataBufferOut(3280) <= dataBufferIn(4016) when (flag_long='1') else '0';
	dataBufferOut(3281) <= dataBufferIn(4759) when (flag_long='1') else '0';
	dataBufferOut(3282) <= dataBufferIn(5502) when (flag_long='1') else '0';
	dataBufferOut(3283) <= dataBufferIn( 101) when (flag_long='1') else '0';
	dataBufferOut(3284) <= dataBufferIn( 844) when (flag_long='1') else '0';
	dataBufferOut(3285) <= dataBufferIn(1587) when (flag_long='1') else '0';
	dataBufferOut(3286) <= dataBufferIn(2330) when (flag_long='1') else '0';
	dataBufferOut(3287) <= dataBufferIn(3073) when (flag_long='1') else '0';
	dataBufferOut(3288) <= dataBufferIn(3816) when (flag_long='1') else '0';
	dataBufferOut(3289) <= dataBufferIn(4559) when (flag_long='1') else '0';
	dataBufferOut(3290) <= dataBufferIn(5302) when (flag_long='1') else '0';
	dataBufferOut(3291) <= dataBufferIn(6045) when (flag_long='1') else '0';
	dataBufferOut(3292) <= dataBufferIn( 644) when (flag_long='1') else '0';
	dataBufferOut(3293) <= dataBufferIn(1387) when (flag_long='1') else '0';
	dataBufferOut(3294) <= dataBufferIn(2130) when (flag_long='1') else '0';
	dataBufferOut(3295) <= dataBufferIn(2873) when (flag_long='1') else '0';
	dataBufferOut(3296) <= dataBufferIn(3616) when (flag_long='1') else '0';
	dataBufferOut(3297) <= dataBufferIn(4359) when (flag_long='1') else '0';
	dataBufferOut(3298) <= dataBufferIn(5102) when (flag_long='1') else '0';
	dataBufferOut(3299) <= dataBufferIn(5845) when (flag_long='1') else '0';
	dataBufferOut(3300) <= dataBufferIn( 444) when (flag_long='1') else '0';
	dataBufferOut(3301) <= dataBufferIn(1187) when (flag_long='1') else '0';
	dataBufferOut(3302) <= dataBufferIn(1930) when (flag_long='1') else '0';
	dataBufferOut(3303) <= dataBufferIn(2673) when (flag_long='1') else '0';
	dataBufferOut(3304) <= dataBufferIn(3416) when (flag_long='1') else '0';
	dataBufferOut(3305) <= dataBufferIn(4159) when (flag_long='1') else '0';
	dataBufferOut(3306) <= dataBufferIn(4902) when (flag_long='1') else '0';
	dataBufferOut(3307) <= dataBufferIn(5645) when (flag_long='1') else '0';
	dataBufferOut(3308) <= dataBufferIn( 244) when (flag_long='1') else '0';
	dataBufferOut(3309) <= dataBufferIn( 987) when (flag_long='1') else '0';
	dataBufferOut(3310) <= dataBufferIn(1730) when (flag_long='1') else '0';
	dataBufferOut(3311) <= dataBufferIn(2473) when (flag_long='1') else '0';
	dataBufferOut(3312) <= dataBufferIn(3216) when (flag_long='1') else '0';
	dataBufferOut(3313) <= dataBufferIn(3959) when (flag_long='1') else '0';
	dataBufferOut(3314) <= dataBufferIn(4702) when (flag_long='1') else '0';
	dataBufferOut(3315) <= dataBufferIn(5445) when (flag_long='1') else '0';
	dataBufferOut(3316) <= dataBufferIn(  44) when (flag_long='1') else '0';
	dataBufferOut(3317) <= dataBufferIn( 787) when (flag_long='1') else '0';
	dataBufferOut(3318) <= dataBufferIn(1530) when (flag_long='1') else '0';
	dataBufferOut(3319) <= dataBufferIn(2273) when (flag_long='1') else '0';
	dataBufferOut(3320) <= dataBufferIn(3016) when (flag_long='1') else '0';
	dataBufferOut(3321) <= dataBufferIn(3759) when (flag_long='1') else '0';
	dataBufferOut(3322) <= dataBufferIn(4502) when (flag_long='1') else '0';
	dataBufferOut(3323) <= dataBufferIn(5245) when (flag_long='1') else '0';
	dataBufferOut(3324) <= dataBufferIn(5988) when (flag_long='1') else '0';
	dataBufferOut(3325) <= dataBufferIn( 587) when (flag_long='1') else '0';
	dataBufferOut(3326) <= dataBufferIn(1330) when (flag_long='1') else '0';
	dataBufferOut(3327) <= dataBufferIn(2073) when (flag_long='1') else '0';
	dataBufferOut(3328) <= dataBufferIn(2816) when (flag_long='1') else '0';
	dataBufferOut(3329) <= dataBufferIn(3559) when (flag_long='1') else '0';
	dataBufferOut(3330) <= dataBufferIn(4302) when (flag_long='1') else '0';
	dataBufferOut(3331) <= dataBufferIn(5045) when (flag_long='1') else '0';
	dataBufferOut(3332) <= dataBufferIn(5788) when (flag_long='1') else '0';
	dataBufferOut(3333) <= dataBufferIn( 387) when (flag_long='1') else '0';
	dataBufferOut(3334) <= dataBufferIn(1130) when (flag_long='1') else '0';
	dataBufferOut(3335) <= dataBufferIn(1873) when (flag_long='1') else '0';
	dataBufferOut(3336) <= dataBufferIn(2616) when (flag_long='1') else '0';
	dataBufferOut(3337) <= dataBufferIn(3359) when (flag_long='1') else '0';
	dataBufferOut(3338) <= dataBufferIn(4102) when (flag_long='1') else '0';
	dataBufferOut(3339) <= dataBufferIn(4845) when (flag_long='1') else '0';
	dataBufferOut(3340) <= dataBufferIn(5588) when (flag_long='1') else '0';
	dataBufferOut(3341) <= dataBufferIn( 187) when (flag_long='1') else '0';
	dataBufferOut(3342) <= dataBufferIn( 930) when (flag_long='1') else '0';
	dataBufferOut(3343) <= dataBufferIn(1673) when (flag_long='1') else '0';
	dataBufferOut(3344) <= dataBufferIn(2416) when (flag_long='1') else '0';
	dataBufferOut(3345) <= dataBufferIn(3159) when (flag_long='1') else '0';
	dataBufferOut(3346) <= dataBufferIn(3902) when (flag_long='1') else '0';
	dataBufferOut(3347) <= dataBufferIn(4645) when (flag_long='1') else '0';
	dataBufferOut(3348) <= dataBufferIn(5388) when (flag_long='1') else '0';
	dataBufferOut(3349) <= dataBufferIn(6131) when (flag_long='1') else '0';
	dataBufferOut(3350) <= dataBufferIn( 730) when (flag_long='1') else '0';
	dataBufferOut(3351) <= dataBufferIn(1473) when (flag_long='1') else '0';
	dataBufferOut(3352) <= dataBufferIn(2216) when (flag_long='1') else '0';
	dataBufferOut(3353) <= dataBufferIn(2959) when (flag_long='1') else '0';
	dataBufferOut(3354) <= dataBufferIn(3702) when (flag_long='1') else '0';
	dataBufferOut(3355) <= dataBufferIn(4445) when (flag_long='1') else '0';
	dataBufferOut(3356) <= dataBufferIn(5188) when (flag_long='1') else '0';
	dataBufferOut(3357) <= dataBufferIn(5931) when (flag_long='1') else '0';
	dataBufferOut(3358) <= dataBufferIn( 530) when (flag_long='1') else '0';
	dataBufferOut(3359) <= dataBufferIn(1273) when (flag_long='1') else '0';
	dataBufferOut(3360) <= dataBufferIn(2016) when (flag_long='1') else '0';
	dataBufferOut(3361) <= dataBufferIn(2759) when (flag_long='1') else '0';
	dataBufferOut(3362) <= dataBufferIn(3502) when (flag_long='1') else '0';
	dataBufferOut(3363) <= dataBufferIn(4245) when (flag_long='1') else '0';
	dataBufferOut(3364) <= dataBufferIn(4988) when (flag_long='1') else '0';
	dataBufferOut(3365) <= dataBufferIn(5731) when (flag_long='1') else '0';
	dataBufferOut(3366) <= dataBufferIn( 330) when (flag_long='1') else '0';
	dataBufferOut(3367) <= dataBufferIn(1073) when (flag_long='1') else '0';
	dataBufferOut(3368) <= dataBufferIn(1816) when (flag_long='1') else '0';
	dataBufferOut(3369) <= dataBufferIn(2559) when (flag_long='1') else '0';
	dataBufferOut(3370) <= dataBufferIn(3302) when (flag_long='1') else '0';
	dataBufferOut(3371) <= dataBufferIn(4045) when (flag_long='1') else '0';
	dataBufferOut(3372) <= dataBufferIn(4788) when (flag_long='1') else '0';
	dataBufferOut(3373) <= dataBufferIn(5531) when (flag_long='1') else '0';
	dataBufferOut(3374) <= dataBufferIn( 130) when (flag_long='1') else '0';
	dataBufferOut(3375) <= dataBufferIn( 873) when (flag_long='1') else '0';
	dataBufferOut(3376) <= dataBufferIn(1616) when (flag_long='1') else '0';
	dataBufferOut(3377) <= dataBufferIn(2359) when (flag_long='1') else '0';
	dataBufferOut(3378) <= dataBufferIn(3102) when (flag_long='1') else '0';
	dataBufferOut(3379) <= dataBufferIn(3845) when (flag_long='1') else '0';
	dataBufferOut(3380) <= dataBufferIn(4588) when (flag_long='1') else '0';
	dataBufferOut(3381) <= dataBufferIn(5331) when (flag_long='1') else '0';
	dataBufferOut(3382) <= dataBufferIn(6074) when (flag_long='1') else '0';
	dataBufferOut(3383) <= dataBufferIn( 673) when (flag_long='1') else '0';
	dataBufferOut(3384) <= dataBufferIn(1416) when (flag_long='1') else '0';
	dataBufferOut(3385) <= dataBufferIn(2159) when (flag_long='1') else '0';
	dataBufferOut(3386) <= dataBufferIn(2902) when (flag_long='1') else '0';
	dataBufferOut(3387) <= dataBufferIn(3645) when (flag_long='1') else '0';
	dataBufferOut(3388) <= dataBufferIn(4388) when (flag_long='1') else '0';
	dataBufferOut(3389) <= dataBufferIn(5131) when (flag_long='1') else '0';
	dataBufferOut(3390) <= dataBufferIn(5874) when (flag_long='1') else '0';
	dataBufferOut(3391) <= dataBufferIn( 473) when (flag_long='1') else '0';
	dataBufferOut(3392) <= dataBufferIn(1216) when (flag_long='1') else '0';
	dataBufferOut(3393) <= dataBufferIn(1959) when (flag_long='1') else '0';
	dataBufferOut(3394) <= dataBufferIn(2702) when (flag_long='1') else '0';
	dataBufferOut(3395) <= dataBufferIn(3445) when (flag_long='1') else '0';
	dataBufferOut(3396) <= dataBufferIn(4188) when (flag_long='1') else '0';
	dataBufferOut(3397) <= dataBufferIn(4931) when (flag_long='1') else '0';
	dataBufferOut(3398) <= dataBufferIn(5674) when (flag_long='1') else '0';
	dataBufferOut(3399) <= dataBufferIn( 273) when (flag_long='1') else '0';
	dataBufferOut(3400) <= dataBufferIn(1016) when (flag_long='1') else '0';
	dataBufferOut(3401) <= dataBufferIn(1759) when (flag_long='1') else '0';
	dataBufferOut(3402) <= dataBufferIn(2502) when (flag_long='1') else '0';
	dataBufferOut(3403) <= dataBufferIn(3245) when (flag_long='1') else '0';
	dataBufferOut(3404) <= dataBufferIn(3988) when (flag_long='1') else '0';
	dataBufferOut(3405) <= dataBufferIn(4731) when (flag_long='1') else '0';
	dataBufferOut(3406) <= dataBufferIn(5474) when (flag_long='1') else '0';
	dataBufferOut(3407) <= dataBufferIn(  73) when (flag_long='1') else '0';
	dataBufferOut(3408) <= dataBufferIn( 816) when (flag_long='1') else '0';
	dataBufferOut(3409) <= dataBufferIn(1559) when (flag_long='1') else '0';
	dataBufferOut(3410) <= dataBufferIn(2302) when (flag_long='1') else '0';
	dataBufferOut(3411) <= dataBufferIn(3045) when (flag_long='1') else '0';
	dataBufferOut(3412) <= dataBufferIn(3788) when (flag_long='1') else '0';
	dataBufferOut(3413) <= dataBufferIn(4531) when (flag_long='1') else '0';
	dataBufferOut(3414) <= dataBufferIn(5274) when (flag_long='1') else '0';
	dataBufferOut(3415) <= dataBufferIn(6017) when (flag_long='1') else '0';
	dataBufferOut(3416) <= dataBufferIn( 616) when (flag_long='1') else '0';
	dataBufferOut(3417) <= dataBufferIn(1359) when (flag_long='1') else '0';
	dataBufferOut(3418) <= dataBufferIn(2102) when (flag_long='1') else '0';
	dataBufferOut(3419) <= dataBufferIn(2845) when (flag_long='1') else '0';
	dataBufferOut(3420) <= dataBufferIn(3588) when (flag_long='1') else '0';
	dataBufferOut(3421) <= dataBufferIn(4331) when (flag_long='1') else '0';
	dataBufferOut(3422) <= dataBufferIn(5074) when (flag_long='1') else '0';
	dataBufferOut(3423) <= dataBufferIn(5817) when (flag_long='1') else '0';
	dataBufferOut(3424) <= dataBufferIn( 416) when (flag_long='1') else '0';
	dataBufferOut(3425) <= dataBufferIn(1159) when (flag_long='1') else '0';
	dataBufferOut(3426) <= dataBufferIn(1902) when (flag_long='1') else '0';
	dataBufferOut(3427) <= dataBufferIn(2645) when (flag_long='1') else '0';
	dataBufferOut(3428) <= dataBufferIn(3388) when (flag_long='1') else '0';
	dataBufferOut(3429) <= dataBufferIn(4131) when (flag_long='1') else '0';
	dataBufferOut(3430) <= dataBufferIn(4874) when (flag_long='1') else '0';
	dataBufferOut(3431) <= dataBufferIn(5617) when (flag_long='1') else '0';
	dataBufferOut(3432) <= dataBufferIn( 216) when (flag_long='1') else '0';
	dataBufferOut(3433) <= dataBufferIn( 959) when (flag_long='1') else '0';
	dataBufferOut(3434) <= dataBufferIn(1702) when (flag_long='1') else '0';
	dataBufferOut(3435) <= dataBufferIn(2445) when (flag_long='1') else '0';
	dataBufferOut(3436) <= dataBufferIn(3188) when (flag_long='1') else '0';
	dataBufferOut(3437) <= dataBufferIn(3931) when (flag_long='1') else '0';
	dataBufferOut(3438) <= dataBufferIn(4674) when (flag_long='1') else '0';
	dataBufferOut(3439) <= dataBufferIn(5417) when (flag_long='1') else '0';
	dataBufferOut(3440) <= dataBufferIn(  16) when (flag_long='1') else '0';
	dataBufferOut(3441) <= dataBufferIn( 759) when (flag_long='1') else '0';
	dataBufferOut(3442) <= dataBufferIn(1502) when (flag_long='1') else '0';
	dataBufferOut(3443) <= dataBufferIn(2245) when (flag_long='1') else '0';
	dataBufferOut(3444) <= dataBufferIn(2988) when (flag_long='1') else '0';
	dataBufferOut(3445) <= dataBufferIn(3731) when (flag_long='1') else '0';
	dataBufferOut(3446) <= dataBufferIn(4474) when (flag_long='1') else '0';
	dataBufferOut(3447) <= dataBufferIn(5217) when (flag_long='1') else '0';
	dataBufferOut(3448) <= dataBufferIn(5960) when (flag_long='1') else '0';
	dataBufferOut(3449) <= dataBufferIn( 559) when (flag_long='1') else '0';
	dataBufferOut(3450) <= dataBufferIn(1302) when (flag_long='1') else '0';
	dataBufferOut(3451) <= dataBufferIn(2045) when (flag_long='1') else '0';
	dataBufferOut(3452) <= dataBufferIn(2788) when (flag_long='1') else '0';
	dataBufferOut(3453) <= dataBufferIn(3531) when (flag_long='1') else '0';
	dataBufferOut(3454) <= dataBufferIn(4274) when (flag_long='1') else '0';
	dataBufferOut(3455) <= dataBufferIn(5017) when (flag_long='1') else '0';
	dataBufferOut(3456) <= dataBufferIn(5760) when (flag_long='1') else '0';
	dataBufferOut(3457) <= dataBufferIn( 359) when (flag_long='1') else '0';
	dataBufferOut(3458) <= dataBufferIn(1102) when (flag_long='1') else '0';
	dataBufferOut(3459) <= dataBufferIn(1845) when (flag_long='1') else '0';
	dataBufferOut(3460) <= dataBufferIn(2588) when (flag_long='1') else '0';
	dataBufferOut(3461) <= dataBufferIn(3331) when (flag_long='1') else '0';
	dataBufferOut(3462) <= dataBufferIn(4074) when (flag_long='1') else '0';
	dataBufferOut(3463) <= dataBufferIn(4817) when (flag_long='1') else '0';
	dataBufferOut(3464) <= dataBufferIn(5560) when (flag_long='1') else '0';
	dataBufferOut(3465) <= dataBufferIn( 159) when (flag_long='1') else '0';
	dataBufferOut(3466) <= dataBufferIn( 902) when (flag_long='1') else '0';
	dataBufferOut(3467) <= dataBufferIn(1645) when (flag_long='1') else '0';
	dataBufferOut(3468) <= dataBufferIn(2388) when (flag_long='1') else '0';
	dataBufferOut(3469) <= dataBufferIn(3131) when (flag_long='1') else '0';
	dataBufferOut(3470) <= dataBufferIn(3874) when (flag_long='1') else '0';
	dataBufferOut(3471) <= dataBufferIn(4617) when (flag_long='1') else '0';
	dataBufferOut(3472) <= dataBufferIn(5360) when (flag_long='1') else '0';
	dataBufferOut(3473) <= dataBufferIn(6103) when (flag_long='1') else '0';
	dataBufferOut(3474) <= dataBufferIn( 702) when (flag_long='1') else '0';
	dataBufferOut(3475) <= dataBufferIn(1445) when (flag_long='1') else '0';
	dataBufferOut(3476) <= dataBufferIn(2188) when (flag_long='1') else '0';
	dataBufferOut(3477) <= dataBufferIn(2931) when (flag_long='1') else '0';
	dataBufferOut(3478) <= dataBufferIn(3674) when (flag_long='1') else '0';
	dataBufferOut(3479) <= dataBufferIn(4417) when (flag_long='1') else '0';
	dataBufferOut(3480) <= dataBufferIn(5160) when (flag_long='1') else '0';
	dataBufferOut(3481) <= dataBufferIn(5903) when (flag_long='1') else '0';
	dataBufferOut(3482) <= dataBufferIn( 502) when (flag_long='1') else '0';
	dataBufferOut(3483) <= dataBufferIn(1245) when (flag_long='1') else '0';
	dataBufferOut(3484) <= dataBufferIn(1988) when (flag_long='1') else '0';
	dataBufferOut(3485) <= dataBufferIn(2731) when (flag_long='1') else '0';
	dataBufferOut(3486) <= dataBufferIn(3474) when (flag_long='1') else '0';
	dataBufferOut(3487) <= dataBufferIn(4217) when (flag_long='1') else '0';
	dataBufferOut(3488) <= dataBufferIn(4960) when (flag_long='1') else '0';
	dataBufferOut(3489) <= dataBufferIn(5703) when (flag_long='1') else '0';
	dataBufferOut(3490) <= dataBufferIn( 302) when (flag_long='1') else '0';
	dataBufferOut(3491) <= dataBufferIn(1045) when (flag_long='1') else '0';
	dataBufferOut(3492) <= dataBufferIn(1788) when (flag_long='1') else '0';
	dataBufferOut(3493) <= dataBufferIn(2531) when (flag_long='1') else '0';
	dataBufferOut(3494) <= dataBufferIn(3274) when (flag_long='1') else '0';
	dataBufferOut(3495) <= dataBufferIn(4017) when (flag_long='1') else '0';
	dataBufferOut(3496) <= dataBufferIn(4760) when (flag_long='1') else '0';
	dataBufferOut(3497) <= dataBufferIn(5503) when (flag_long='1') else '0';
	dataBufferOut(3498) <= dataBufferIn( 102) when (flag_long='1') else '0';
	dataBufferOut(3499) <= dataBufferIn( 845) when (flag_long='1') else '0';
	dataBufferOut(3500) <= dataBufferIn(1588) when (flag_long='1') else '0';
	dataBufferOut(3501) <= dataBufferIn(2331) when (flag_long='1') else '0';
	dataBufferOut(3502) <= dataBufferIn(3074) when (flag_long='1') else '0';
	dataBufferOut(3503) <= dataBufferIn(3817) when (flag_long='1') else '0';
	dataBufferOut(3504) <= dataBufferIn(4560) when (flag_long='1') else '0';
	dataBufferOut(3505) <= dataBufferIn(5303) when (flag_long='1') else '0';
	dataBufferOut(3506) <= dataBufferIn(6046) when (flag_long='1') else '0';
	dataBufferOut(3507) <= dataBufferIn( 645) when (flag_long='1') else '0';
	dataBufferOut(3508) <= dataBufferIn(1388) when (flag_long='1') else '0';
	dataBufferOut(3509) <= dataBufferIn(2131) when (flag_long='1') else '0';
	dataBufferOut(3510) <= dataBufferIn(2874) when (flag_long='1') else '0';
	dataBufferOut(3511) <= dataBufferIn(3617) when (flag_long='1') else '0';
	dataBufferOut(3512) <= dataBufferIn(4360) when (flag_long='1') else '0';
	dataBufferOut(3513) <= dataBufferIn(5103) when (flag_long='1') else '0';
	dataBufferOut(3514) <= dataBufferIn(5846) when (flag_long='1') else '0';
	dataBufferOut(3515) <= dataBufferIn( 445) when (flag_long='1') else '0';
	dataBufferOut(3516) <= dataBufferIn(1188) when (flag_long='1') else '0';
	dataBufferOut(3517) <= dataBufferIn(1931) when (flag_long='1') else '0';
	dataBufferOut(3518) <= dataBufferIn(2674) when (flag_long='1') else '0';
	dataBufferOut(3519) <= dataBufferIn(3417) when (flag_long='1') else '0';
	dataBufferOut(3520) <= dataBufferIn(4160) when (flag_long='1') else '0';
	dataBufferOut(3521) <= dataBufferIn(4903) when (flag_long='1') else '0';
	dataBufferOut(3522) <= dataBufferIn(5646) when (flag_long='1') else '0';
	dataBufferOut(3523) <= dataBufferIn( 245) when (flag_long='1') else '0';
	dataBufferOut(3524) <= dataBufferIn( 988) when (flag_long='1') else '0';
	dataBufferOut(3525) <= dataBufferIn(1731) when (flag_long='1') else '0';
	dataBufferOut(3526) <= dataBufferIn(2474) when (flag_long='1') else '0';
	dataBufferOut(3527) <= dataBufferIn(3217) when (flag_long='1') else '0';
	dataBufferOut(3528) <= dataBufferIn(3960) when (flag_long='1') else '0';
	dataBufferOut(3529) <= dataBufferIn(4703) when (flag_long='1') else '0';
	dataBufferOut(3530) <= dataBufferIn(5446) when (flag_long='1') else '0';
	dataBufferOut(3531) <= dataBufferIn(  45) when (flag_long='1') else '0';
	dataBufferOut(3532) <= dataBufferIn( 788) when (flag_long='1') else '0';
	dataBufferOut(3533) <= dataBufferIn(1531) when (flag_long='1') else '0';
	dataBufferOut(3534) <= dataBufferIn(2274) when (flag_long='1') else '0';
	dataBufferOut(3535) <= dataBufferIn(3017) when (flag_long='1') else '0';
	dataBufferOut(3536) <= dataBufferIn(3760) when (flag_long='1') else '0';
	dataBufferOut(3537) <= dataBufferIn(4503) when (flag_long='1') else '0';
	dataBufferOut(3538) <= dataBufferIn(5246) when (flag_long='1') else '0';
	dataBufferOut(3539) <= dataBufferIn(5989) when (flag_long='1') else '0';
	dataBufferOut(3540) <= dataBufferIn( 588) when (flag_long='1') else '0';
	dataBufferOut(3541) <= dataBufferIn(1331) when (flag_long='1') else '0';
	dataBufferOut(3542) <= dataBufferIn(2074) when (flag_long='1') else '0';
	dataBufferOut(3543) <= dataBufferIn(2817) when (flag_long='1') else '0';
	dataBufferOut(3544) <= dataBufferIn(3560) when (flag_long='1') else '0';
	dataBufferOut(3545) <= dataBufferIn(4303) when (flag_long='1') else '0';
	dataBufferOut(3546) <= dataBufferIn(5046) when (flag_long='1') else '0';
	dataBufferOut(3547) <= dataBufferIn(5789) when (flag_long='1') else '0';
	dataBufferOut(3548) <= dataBufferIn( 388) when (flag_long='1') else '0';
	dataBufferOut(3549) <= dataBufferIn(1131) when (flag_long='1') else '0';
	dataBufferOut(3550) <= dataBufferIn(1874) when (flag_long='1') else '0';
	dataBufferOut(3551) <= dataBufferIn(2617) when (flag_long='1') else '0';
	dataBufferOut(3552) <= dataBufferIn(3360) when (flag_long='1') else '0';
	dataBufferOut(3553) <= dataBufferIn(4103) when (flag_long='1') else '0';
	dataBufferOut(3554) <= dataBufferIn(4846) when (flag_long='1') else '0';
	dataBufferOut(3555) <= dataBufferIn(5589) when (flag_long='1') else '0';
	dataBufferOut(3556) <= dataBufferIn( 188) when (flag_long='1') else '0';
	dataBufferOut(3557) <= dataBufferIn( 931) when (flag_long='1') else '0';
	dataBufferOut(3558) <= dataBufferIn(1674) when (flag_long='1') else '0';
	dataBufferOut(3559) <= dataBufferIn(2417) when (flag_long='1') else '0';
	dataBufferOut(3560) <= dataBufferIn(3160) when (flag_long='1') else '0';
	dataBufferOut(3561) <= dataBufferIn(3903) when (flag_long='1') else '0';
	dataBufferOut(3562) <= dataBufferIn(4646) when (flag_long='1') else '0';
	dataBufferOut(3563) <= dataBufferIn(5389) when (flag_long='1') else '0';
	dataBufferOut(3564) <= dataBufferIn(6132) when (flag_long='1') else '0';
	dataBufferOut(3565) <= dataBufferIn( 731) when (flag_long='1') else '0';
	dataBufferOut(3566) <= dataBufferIn(1474) when (flag_long='1') else '0';
	dataBufferOut(3567) <= dataBufferIn(2217) when (flag_long='1') else '0';
	dataBufferOut(3568) <= dataBufferIn(2960) when (flag_long='1') else '0';
	dataBufferOut(3569) <= dataBufferIn(3703) when (flag_long='1') else '0';
	dataBufferOut(3570) <= dataBufferIn(4446) when (flag_long='1') else '0';
	dataBufferOut(3571) <= dataBufferIn(5189) when (flag_long='1') else '0';
	dataBufferOut(3572) <= dataBufferIn(5932) when (flag_long='1') else '0';
	dataBufferOut(3573) <= dataBufferIn( 531) when (flag_long='1') else '0';
	dataBufferOut(3574) <= dataBufferIn(1274) when (flag_long='1') else '0';
	dataBufferOut(3575) <= dataBufferIn(2017) when (flag_long='1') else '0';
	dataBufferOut(3576) <= dataBufferIn(2760) when (flag_long='1') else '0';
	dataBufferOut(3577) <= dataBufferIn(3503) when (flag_long='1') else '0';
	dataBufferOut(3578) <= dataBufferIn(4246) when (flag_long='1') else '0';
	dataBufferOut(3579) <= dataBufferIn(4989) when (flag_long='1') else '0';
	dataBufferOut(3580) <= dataBufferIn(5732) when (flag_long='1') else '0';
	dataBufferOut(3581) <= dataBufferIn( 331) when (flag_long='1') else '0';
	dataBufferOut(3582) <= dataBufferIn(1074) when (flag_long='1') else '0';
	dataBufferOut(3583) <= dataBufferIn(1817) when (flag_long='1') else '0';
	dataBufferOut(3584) <= dataBufferIn(2560) when (flag_long='1') else '0';
	dataBufferOut(3585) <= dataBufferIn(3303) when (flag_long='1') else '0';
	dataBufferOut(3586) <= dataBufferIn(4046) when (flag_long='1') else '0';
	dataBufferOut(3587) <= dataBufferIn(4789) when (flag_long='1') else '0';
	dataBufferOut(3588) <= dataBufferIn(5532) when (flag_long='1') else '0';
	dataBufferOut(3589) <= dataBufferIn( 131) when (flag_long='1') else '0';
	dataBufferOut(3590) <= dataBufferIn( 874) when (flag_long='1') else '0';
	dataBufferOut(3591) <= dataBufferIn(1617) when (flag_long='1') else '0';
	dataBufferOut(3592) <= dataBufferIn(2360) when (flag_long='1') else '0';
	dataBufferOut(3593) <= dataBufferIn(3103) when (flag_long='1') else '0';
	dataBufferOut(3594) <= dataBufferIn(3846) when (flag_long='1') else '0';
	dataBufferOut(3595) <= dataBufferIn(4589) when (flag_long='1') else '0';
	dataBufferOut(3596) <= dataBufferIn(5332) when (flag_long='1') else '0';
	dataBufferOut(3597) <= dataBufferIn(6075) when (flag_long='1') else '0';
	dataBufferOut(3598) <= dataBufferIn( 674) when (flag_long='1') else '0';
	dataBufferOut(3599) <= dataBufferIn(1417) when (flag_long='1') else '0';
	dataBufferOut(3600) <= dataBufferIn(2160) when (flag_long='1') else '0';
	dataBufferOut(3601) <= dataBufferIn(2903) when (flag_long='1') else '0';
	dataBufferOut(3602) <= dataBufferIn(3646) when (flag_long='1') else '0';
	dataBufferOut(3603) <= dataBufferIn(4389) when (flag_long='1') else '0';
	dataBufferOut(3604) <= dataBufferIn(5132) when (flag_long='1') else '0';
	dataBufferOut(3605) <= dataBufferIn(5875) when (flag_long='1') else '0';
	dataBufferOut(3606) <= dataBufferIn( 474) when (flag_long='1') else '0';
	dataBufferOut(3607) <= dataBufferIn(1217) when (flag_long='1') else '0';
	dataBufferOut(3608) <= dataBufferIn(1960) when (flag_long='1') else '0';
	dataBufferOut(3609) <= dataBufferIn(2703) when (flag_long='1') else '0';
	dataBufferOut(3610) <= dataBufferIn(3446) when (flag_long='1') else '0';
	dataBufferOut(3611) <= dataBufferIn(4189) when (flag_long='1') else '0';
	dataBufferOut(3612) <= dataBufferIn(4932) when (flag_long='1') else '0';
	dataBufferOut(3613) <= dataBufferIn(5675) when (flag_long='1') else '0';
	dataBufferOut(3614) <= dataBufferIn( 274) when (flag_long='1') else '0';
	dataBufferOut(3615) <= dataBufferIn(1017) when (flag_long='1') else '0';
	dataBufferOut(3616) <= dataBufferIn(1760) when (flag_long='1') else '0';
	dataBufferOut(3617) <= dataBufferIn(2503) when (flag_long='1') else '0';
	dataBufferOut(3618) <= dataBufferIn(3246) when (flag_long='1') else '0';
	dataBufferOut(3619) <= dataBufferIn(3989) when (flag_long='1') else '0';
	dataBufferOut(3620) <= dataBufferIn(4732) when (flag_long='1') else '0';
	dataBufferOut(3621) <= dataBufferIn(5475) when (flag_long='1') else '0';
	dataBufferOut(3622) <= dataBufferIn(  74) when (flag_long='1') else '0';
	dataBufferOut(3623) <= dataBufferIn( 817) when (flag_long='1') else '0';
	dataBufferOut(3624) <= dataBufferIn(1560) when (flag_long='1') else '0';
	dataBufferOut(3625) <= dataBufferIn(2303) when (flag_long='1') else '0';
	dataBufferOut(3626) <= dataBufferIn(3046) when (flag_long='1') else '0';
	dataBufferOut(3627) <= dataBufferIn(3789) when (flag_long='1') else '0';
	dataBufferOut(3628) <= dataBufferIn(4532) when (flag_long='1') else '0';
	dataBufferOut(3629) <= dataBufferIn(5275) when (flag_long='1') else '0';
	dataBufferOut(3630) <= dataBufferIn(6018) when (flag_long='1') else '0';
	dataBufferOut(3631) <= dataBufferIn( 617) when (flag_long='1') else '0';
	dataBufferOut(3632) <= dataBufferIn(1360) when (flag_long='1') else '0';
	dataBufferOut(3633) <= dataBufferIn(2103) when (flag_long='1') else '0';
	dataBufferOut(3634) <= dataBufferIn(2846) when (flag_long='1') else '0';
	dataBufferOut(3635) <= dataBufferIn(3589) when (flag_long='1') else '0';
	dataBufferOut(3636) <= dataBufferIn(4332) when (flag_long='1') else '0';
	dataBufferOut(3637) <= dataBufferIn(5075) when (flag_long='1') else '0';
	dataBufferOut(3638) <= dataBufferIn(5818) when (flag_long='1') else '0';
	dataBufferOut(3639) <= dataBufferIn( 417) when (flag_long='1') else '0';
	dataBufferOut(3640) <= dataBufferIn(1160) when (flag_long='1') else '0';
	dataBufferOut(3641) <= dataBufferIn(1903) when (flag_long='1') else '0';
	dataBufferOut(3642) <= dataBufferIn(2646) when (flag_long='1') else '0';
	dataBufferOut(3643) <= dataBufferIn(3389) when (flag_long='1') else '0';
	dataBufferOut(3644) <= dataBufferIn(4132) when (flag_long='1') else '0';
	dataBufferOut(3645) <= dataBufferIn(4875) when (flag_long='1') else '0';
	dataBufferOut(3646) <= dataBufferIn(5618) when (flag_long='1') else '0';
	dataBufferOut(3647) <= dataBufferIn( 217) when (flag_long='1') else '0';
	dataBufferOut(3648) <= dataBufferIn( 960) when (flag_long='1') else '0';
	dataBufferOut(3649) <= dataBufferIn(1703) when (flag_long='1') else '0';
	dataBufferOut(3650) <= dataBufferIn(2446) when (flag_long='1') else '0';
	dataBufferOut(3651) <= dataBufferIn(3189) when (flag_long='1') else '0';
	dataBufferOut(3652) <= dataBufferIn(3932) when (flag_long='1') else '0';
	dataBufferOut(3653) <= dataBufferIn(4675) when (flag_long='1') else '0';
	dataBufferOut(3654) <= dataBufferIn(5418) when (flag_long='1') else '0';
	dataBufferOut(3655) <= dataBufferIn(  17) when (flag_long='1') else '0';
	dataBufferOut(3656) <= dataBufferIn( 760) when (flag_long='1') else '0';
	dataBufferOut(3657) <= dataBufferIn(1503) when (flag_long='1') else '0';
	dataBufferOut(3658) <= dataBufferIn(2246) when (flag_long='1') else '0';
	dataBufferOut(3659) <= dataBufferIn(2989) when (flag_long='1') else '0';
	dataBufferOut(3660) <= dataBufferIn(3732) when (flag_long='1') else '0';
	dataBufferOut(3661) <= dataBufferIn(4475) when (flag_long='1') else '0';
	dataBufferOut(3662) <= dataBufferIn(5218) when (flag_long='1') else '0';
	dataBufferOut(3663) <= dataBufferIn(5961) when (flag_long='1') else '0';
	dataBufferOut(3664) <= dataBufferIn( 560) when (flag_long='1') else '0';
	dataBufferOut(3665) <= dataBufferIn(1303) when (flag_long='1') else '0';
	dataBufferOut(3666) <= dataBufferIn(2046) when (flag_long='1') else '0';
	dataBufferOut(3667) <= dataBufferIn(2789) when (flag_long='1') else '0';
	dataBufferOut(3668) <= dataBufferIn(3532) when (flag_long='1') else '0';
	dataBufferOut(3669) <= dataBufferIn(4275) when (flag_long='1') else '0';
	dataBufferOut(3670) <= dataBufferIn(5018) when (flag_long='1') else '0';
	dataBufferOut(3671) <= dataBufferIn(5761) when (flag_long='1') else '0';
	dataBufferOut(3672) <= dataBufferIn( 360) when (flag_long='1') else '0';
	dataBufferOut(3673) <= dataBufferIn(1103) when (flag_long='1') else '0';
	dataBufferOut(3674) <= dataBufferIn(1846) when (flag_long='1') else '0';
	dataBufferOut(3675) <= dataBufferIn(2589) when (flag_long='1') else '0';
	dataBufferOut(3676) <= dataBufferIn(3332) when (flag_long='1') else '0';
	dataBufferOut(3677) <= dataBufferIn(4075) when (flag_long='1') else '0';
	dataBufferOut(3678) <= dataBufferIn(4818) when (flag_long='1') else '0';
	dataBufferOut(3679) <= dataBufferIn(5561) when (flag_long='1') else '0';
	dataBufferOut(3680) <= dataBufferIn( 160) when (flag_long='1') else '0';
	dataBufferOut(3681) <= dataBufferIn( 903) when (flag_long='1') else '0';
	dataBufferOut(3682) <= dataBufferIn(1646) when (flag_long='1') else '0';
	dataBufferOut(3683) <= dataBufferIn(2389) when (flag_long='1') else '0';
	dataBufferOut(3684) <= dataBufferIn(3132) when (flag_long='1') else '0';
	dataBufferOut(3685) <= dataBufferIn(3875) when (flag_long='1') else '0';
	dataBufferOut(3686) <= dataBufferIn(4618) when (flag_long='1') else '0';
	dataBufferOut(3687) <= dataBufferIn(5361) when (flag_long='1') else '0';
	dataBufferOut(3688) <= dataBufferIn(6104) when (flag_long='1') else '0';
	dataBufferOut(3689) <= dataBufferIn( 703) when (flag_long='1') else '0';
	dataBufferOut(3690) <= dataBufferIn(1446) when (flag_long='1') else '0';
	dataBufferOut(3691) <= dataBufferIn(2189) when (flag_long='1') else '0';
	dataBufferOut(3692) <= dataBufferIn(2932) when (flag_long='1') else '0';
	dataBufferOut(3693) <= dataBufferIn(3675) when (flag_long='1') else '0';
	dataBufferOut(3694) <= dataBufferIn(4418) when (flag_long='1') else '0';
	dataBufferOut(3695) <= dataBufferIn(5161) when (flag_long='1') else '0';
	dataBufferOut(3696) <= dataBufferIn(5904) when (flag_long='1') else '0';
	dataBufferOut(3697) <= dataBufferIn( 503) when (flag_long='1') else '0';
	dataBufferOut(3698) <= dataBufferIn(1246) when (flag_long='1') else '0';
	dataBufferOut(3699) <= dataBufferIn(1989) when (flag_long='1') else '0';
	dataBufferOut(3700) <= dataBufferIn(2732) when (flag_long='1') else '0';
	dataBufferOut(3701) <= dataBufferIn(3475) when (flag_long='1') else '0';
	dataBufferOut(3702) <= dataBufferIn(4218) when (flag_long='1') else '0';
	dataBufferOut(3703) <= dataBufferIn(4961) when (flag_long='1') else '0';
	dataBufferOut(3704) <= dataBufferIn(5704) when (flag_long='1') else '0';
	dataBufferOut(3705) <= dataBufferIn( 303) when (flag_long='1') else '0';
	dataBufferOut(3706) <= dataBufferIn(1046) when (flag_long='1') else '0';
	dataBufferOut(3707) <= dataBufferIn(1789) when (flag_long='1') else '0';
	dataBufferOut(3708) <= dataBufferIn(2532) when (flag_long='1') else '0';
	dataBufferOut(3709) <= dataBufferIn(3275) when (flag_long='1') else '0';
	dataBufferOut(3710) <= dataBufferIn(4018) when (flag_long='1') else '0';
	dataBufferOut(3711) <= dataBufferIn(4761) when (flag_long='1') else '0';
	dataBufferOut(3712) <= dataBufferIn(5504) when (flag_long='1') else '0';
	dataBufferOut(3713) <= dataBufferIn( 103) when (flag_long='1') else '0';
	dataBufferOut(3714) <= dataBufferIn( 846) when (flag_long='1') else '0';
	dataBufferOut(3715) <= dataBufferIn(1589) when (flag_long='1') else '0';
	dataBufferOut(3716) <= dataBufferIn(2332) when (flag_long='1') else '0';
	dataBufferOut(3717) <= dataBufferIn(3075) when (flag_long='1') else '0';
	dataBufferOut(3718) <= dataBufferIn(3818) when (flag_long='1') else '0';
	dataBufferOut(3719) <= dataBufferIn(4561) when (flag_long='1') else '0';
	dataBufferOut(3720) <= dataBufferIn(5304) when (flag_long='1') else '0';
	dataBufferOut(3721) <= dataBufferIn(6047) when (flag_long='1') else '0';
	dataBufferOut(3722) <= dataBufferIn( 646) when (flag_long='1') else '0';
	dataBufferOut(3723) <= dataBufferIn(1389) when (flag_long='1') else '0';
	dataBufferOut(3724) <= dataBufferIn(2132) when (flag_long='1') else '0';
	dataBufferOut(3725) <= dataBufferIn(2875) when (flag_long='1') else '0';
	dataBufferOut(3726) <= dataBufferIn(3618) when (flag_long='1') else '0';
	dataBufferOut(3727) <= dataBufferIn(4361) when (flag_long='1') else '0';
	dataBufferOut(3728) <= dataBufferIn(5104) when (flag_long='1') else '0';
	dataBufferOut(3729) <= dataBufferIn(5847) when (flag_long='1') else '0';
	dataBufferOut(3730) <= dataBufferIn( 446) when (flag_long='1') else '0';
	dataBufferOut(3731) <= dataBufferIn(1189) when (flag_long='1') else '0';
	dataBufferOut(3732) <= dataBufferIn(1932) when (flag_long='1') else '0';
	dataBufferOut(3733) <= dataBufferIn(2675) when (flag_long='1') else '0';
	dataBufferOut(3734) <= dataBufferIn(3418) when (flag_long='1') else '0';
	dataBufferOut(3735) <= dataBufferIn(4161) when (flag_long='1') else '0';
	dataBufferOut(3736) <= dataBufferIn(4904) when (flag_long='1') else '0';
	dataBufferOut(3737) <= dataBufferIn(5647) when (flag_long='1') else '0';
	dataBufferOut(3738) <= dataBufferIn( 246) when (flag_long='1') else '0';
	dataBufferOut(3739) <= dataBufferIn( 989) when (flag_long='1') else '0';
	dataBufferOut(3740) <= dataBufferIn(1732) when (flag_long='1') else '0';
	dataBufferOut(3741) <= dataBufferIn(2475) when (flag_long='1') else '0';
	dataBufferOut(3742) <= dataBufferIn(3218) when (flag_long='1') else '0';
	dataBufferOut(3743) <= dataBufferIn(3961) when (flag_long='1') else '0';
	dataBufferOut(3744) <= dataBufferIn(4704) when (flag_long='1') else '0';
	dataBufferOut(3745) <= dataBufferIn(5447) when (flag_long='1') else '0';
	dataBufferOut(3746) <= dataBufferIn(  46) when (flag_long='1') else '0';
	dataBufferOut(3747) <= dataBufferIn( 789) when (flag_long='1') else '0';
	dataBufferOut(3748) <= dataBufferIn(1532) when (flag_long='1') else '0';
	dataBufferOut(3749) <= dataBufferIn(2275) when (flag_long='1') else '0';
	dataBufferOut(3750) <= dataBufferIn(3018) when (flag_long='1') else '0';
	dataBufferOut(3751) <= dataBufferIn(3761) when (flag_long='1') else '0';
	dataBufferOut(3752) <= dataBufferIn(4504) when (flag_long='1') else '0';
	dataBufferOut(3753) <= dataBufferIn(5247) when (flag_long='1') else '0';
	dataBufferOut(3754) <= dataBufferIn(5990) when (flag_long='1') else '0';
	dataBufferOut(3755) <= dataBufferIn( 589) when (flag_long='1') else '0';
	dataBufferOut(3756) <= dataBufferIn(1332) when (flag_long='1') else '0';
	dataBufferOut(3757) <= dataBufferIn(2075) when (flag_long='1') else '0';
	dataBufferOut(3758) <= dataBufferIn(2818) when (flag_long='1') else '0';
	dataBufferOut(3759) <= dataBufferIn(3561) when (flag_long='1') else '0';
	dataBufferOut(3760) <= dataBufferIn(4304) when (flag_long='1') else '0';
	dataBufferOut(3761) <= dataBufferIn(5047) when (flag_long='1') else '0';
	dataBufferOut(3762) <= dataBufferIn(5790) when (flag_long='1') else '0';
	dataBufferOut(3763) <= dataBufferIn( 389) when (flag_long='1') else '0';
	dataBufferOut(3764) <= dataBufferIn(1132) when (flag_long='1') else '0';
	dataBufferOut(3765) <= dataBufferIn(1875) when (flag_long='1') else '0';
	dataBufferOut(3766) <= dataBufferIn(2618) when (flag_long='1') else '0';
	dataBufferOut(3767) <= dataBufferIn(3361) when (flag_long='1') else '0';
	dataBufferOut(3768) <= dataBufferIn(4104) when (flag_long='1') else '0';
	dataBufferOut(3769) <= dataBufferIn(4847) when (flag_long='1') else '0';
	dataBufferOut(3770) <= dataBufferIn(5590) when (flag_long='1') else '0';
	dataBufferOut(3771) <= dataBufferIn( 189) when (flag_long='1') else '0';
	dataBufferOut(3772) <= dataBufferIn( 932) when (flag_long='1') else '0';
	dataBufferOut(3773) <= dataBufferIn(1675) when (flag_long='1') else '0';
	dataBufferOut(3774) <= dataBufferIn(2418) when (flag_long='1') else '0';
	dataBufferOut(3775) <= dataBufferIn(3161) when (flag_long='1') else '0';
	dataBufferOut(3776) <= dataBufferIn(3904) when (flag_long='1') else '0';
	dataBufferOut(3777) <= dataBufferIn(4647) when (flag_long='1') else '0';
	dataBufferOut(3778) <= dataBufferIn(5390) when (flag_long='1') else '0';
	dataBufferOut(3779) <= dataBufferIn(6133) when (flag_long='1') else '0';
	dataBufferOut(3780) <= dataBufferIn( 732) when (flag_long='1') else '0';
	dataBufferOut(3781) <= dataBufferIn(1475) when (flag_long='1') else '0';
	dataBufferOut(3782) <= dataBufferIn(2218) when (flag_long='1') else '0';
	dataBufferOut(3783) <= dataBufferIn(2961) when (flag_long='1') else '0';
	dataBufferOut(3784) <= dataBufferIn(3704) when (flag_long='1') else '0';
	dataBufferOut(3785) <= dataBufferIn(4447) when (flag_long='1') else '0';
	dataBufferOut(3786) <= dataBufferIn(5190) when (flag_long='1') else '0';
	dataBufferOut(3787) <= dataBufferIn(5933) when (flag_long='1') else '0';
	dataBufferOut(3788) <= dataBufferIn( 532) when (flag_long='1') else '0';
	dataBufferOut(3789) <= dataBufferIn(1275) when (flag_long='1') else '0';
	dataBufferOut(3790) <= dataBufferIn(2018) when (flag_long='1') else '0';
	dataBufferOut(3791) <= dataBufferIn(2761) when (flag_long='1') else '0';
	dataBufferOut(3792) <= dataBufferIn(3504) when (flag_long='1') else '0';
	dataBufferOut(3793) <= dataBufferIn(4247) when (flag_long='1') else '0';
	dataBufferOut(3794) <= dataBufferIn(4990) when (flag_long='1') else '0';
	dataBufferOut(3795) <= dataBufferIn(5733) when (flag_long='1') else '0';
	dataBufferOut(3796) <= dataBufferIn( 332) when (flag_long='1') else '0';
	dataBufferOut(3797) <= dataBufferIn(1075) when (flag_long='1') else '0';
	dataBufferOut(3798) <= dataBufferIn(1818) when (flag_long='1') else '0';
	dataBufferOut(3799) <= dataBufferIn(2561) when (flag_long='1') else '0';
	dataBufferOut(3800) <= dataBufferIn(3304) when (flag_long='1') else '0';
	dataBufferOut(3801) <= dataBufferIn(4047) when (flag_long='1') else '0';
	dataBufferOut(3802) <= dataBufferIn(4790) when (flag_long='1') else '0';
	dataBufferOut(3803) <= dataBufferIn(5533) when (flag_long='1') else '0';
	dataBufferOut(3804) <= dataBufferIn( 132) when (flag_long='1') else '0';
	dataBufferOut(3805) <= dataBufferIn( 875) when (flag_long='1') else '0';
	dataBufferOut(3806) <= dataBufferIn(1618) when (flag_long='1') else '0';
	dataBufferOut(3807) <= dataBufferIn(2361) when (flag_long='1') else '0';
	dataBufferOut(3808) <= dataBufferIn(3104) when (flag_long='1') else '0';
	dataBufferOut(3809) <= dataBufferIn(3847) when (flag_long='1') else '0';
	dataBufferOut(3810) <= dataBufferIn(4590) when (flag_long='1') else '0';
	dataBufferOut(3811) <= dataBufferIn(5333) when (flag_long='1') else '0';
	dataBufferOut(3812) <= dataBufferIn(6076) when (flag_long='1') else '0';
	dataBufferOut(3813) <= dataBufferIn( 675) when (flag_long='1') else '0';
	dataBufferOut(3814) <= dataBufferIn(1418) when (flag_long='1') else '0';
	dataBufferOut(3815) <= dataBufferIn(2161) when (flag_long='1') else '0';
	dataBufferOut(3816) <= dataBufferIn(2904) when (flag_long='1') else '0';
	dataBufferOut(3817) <= dataBufferIn(3647) when (flag_long='1') else '0';
	dataBufferOut(3818) <= dataBufferIn(4390) when (flag_long='1') else '0';
	dataBufferOut(3819) <= dataBufferIn(5133) when (flag_long='1') else '0';
	dataBufferOut(3820) <= dataBufferIn(5876) when (flag_long='1') else '0';
	dataBufferOut(3821) <= dataBufferIn( 475) when (flag_long='1') else '0';
	dataBufferOut(3822) <= dataBufferIn(1218) when (flag_long='1') else '0';
	dataBufferOut(3823) <= dataBufferIn(1961) when (flag_long='1') else '0';
	dataBufferOut(3824) <= dataBufferIn(2704) when (flag_long='1') else '0';
	dataBufferOut(3825) <= dataBufferIn(3447) when (flag_long='1') else '0';
	dataBufferOut(3826) <= dataBufferIn(4190) when (flag_long='1') else '0';
	dataBufferOut(3827) <= dataBufferIn(4933) when (flag_long='1') else '0';
	dataBufferOut(3828) <= dataBufferIn(5676) when (flag_long='1') else '0';
	dataBufferOut(3829) <= dataBufferIn( 275) when (flag_long='1') else '0';
	dataBufferOut(3830) <= dataBufferIn(1018) when (flag_long='1') else '0';
	dataBufferOut(3831) <= dataBufferIn(1761) when (flag_long='1') else '0';
	dataBufferOut(3832) <= dataBufferIn(2504) when (flag_long='1') else '0';
	dataBufferOut(3833) <= dataBufferIn(3247) when (flag_long='1') else '0';
	dataBufferOut(3834) <= dataBufferIn(3990) when (flag_long='1') else '0';
	dataBufferOut(3835) <= dataBufferIn(4733) when (flag_long='1') else '0';
	dataBufferOut(3836) <= dataBufferIn(5476) when (flag_long='1') else '0';
	dataBufferOut(3837) <= dataBufferIn(  75) when (flag_long='1') else '0';
	dataBufferOut(3838) <= dataBufferIn( 818) when (flag_long='1') else '0';
	dataBufferOut(3839) <= dataBufferIn(1561) when (flag_long='1') else '0';
	dataBufferOut(3840) <= dataBufferIn(2304) when (flag_long='1') else '0';
	dataBufferOut(3841) <= dataBufferIn(3047) when (flag_long='1') else '0';
	dataBufferOut(3842) <= dataBufferIn(3790) when (flag_long='1') else '0';
	dataBufferOut(3843) <= dataBufferIn(4533) when (flag_long='1') else '0';
	dataBufferOut(3844) <= dataBufferIn(5276) when (flag_long='1') else '0';
	dataBufferOut(3845) <= dataBufferIn(6019) when (flag_long='1') else '0';
	dataBufferOut(3846) <= dataBufferIn( 618) when (flag_long='1') else '0';
	dataBufferOut(3847) <= dataBufferIn(1361) when (flag_long='1') else '0';
	dataBufferOut(3848) <= dataBufferIn(2104) when (flag_long='1') else '0';
	dataBufferOut(3849) <= dataBufferIn(2847) when (flag_long='1') else '0';
	dataBufferOut(3850) <= dataBufferIn(3590) when (flag_long='1') else '0';
	dataBufferOut(3851) <= dataBufferIn(4333) when (flag_long='1') else '0';
	dataBufferOut(3852) <= dataBufferIn(5076) when (flag_long='1') else '0';
	dataBufferOut(3853) <= dataBufferIn(5819) when (flag_long='1') else '0';
	dataBufferOut(3854) <= dataBufferIn( 418) when (flag_long='1') else '0';
	dataBufferOut(3855) <= dataBufferIn(1161) when (flag_long='1') else '0';
	dataBufferOut(3856) <= dataBufferIn(1904) when (flag_long='1') else '0';
	dataBufferOut(3857) <= dataBufferIn(2647) when (flag_long='1') else '0';
	dataBufferOut(3858) <= dataBufferIn(3390) when (flag_long='1') else '0';
	dataBufferOut(3859) <= dataBufferIn(4133) when (flag_long='1') else '0';
	dataBufferOut(3860) <= dataBufferIn(4876) when (flag_long='1') else '0';
	dataBufferOut(3861) <= dataBufferIn(5619) when (flag_long='1') else '0';
	dataBufferOut(3862) <= dataBufferIn( 218) when (flag_long='1') else '0';
	dataBufferOut(3863) <= dataBufferIn( 961) when (flag_long='1') else '0';
	dataBufferOut(3864) <= dataBufferIn(1704) when (flag_long='1') else '0';
	dataBufferOut(3865) <= dataBufferIn(2447) when (flag_long='1') else '0';
	dataBufferOut(3866) <= dataBufferIn(3190) when (flag_long='1') else '0';
	dataBufferOut(3867) <= dataBufferIn(3933) when (flag_long='1') else '0';
	dataBufferOut(3868) <= dataBufferIn(4676) when (flag_long='1') else '0';
	dataBufferOut(3869) <= dataBufferIn(5419) when (flag_long='1') else '0';
	dataBufferOut(3870) <= dataBufferIn(  18) when (flag_long='1') else '0';
	dataBufferOut(3871) <= dataBufferIn( 761) when (flag_long='1') else '0';
	dataBufferOut(3872) <= dataBufferIn(1504) when (flag_long='1') else '0';
	dataBufferOut(3873) <= dataBufferIn(2247) when (flag_long='1') else '0';
	dataBufferOut(3874) <= dataBufferIn(2990) when (flag_long='1') else '0';
	dataBufferOut(3875) <= dataBufferIn(3733) when (flag_long='1') else '0';
	dataBufferOut(3876) <= dataBufferIn(4476) when (flag_long='1') else '0';
	dataBufferOut(3877) <= dataBufferIn(5219) when (flag_long='1') else '0';
	dataBufferOut(3878) <= dataBufferIn(5962) when (flag_long='1') else '0';
	dataBufferOut(3879) <= dataBufferIn( 561) when (flag_long='1') else '0';
	dataBufferOut(3880) <= dataBufferIn(1304) when (flag_long='1') else '0';
	dataBufferOut(3881) <= dataBufferIn(2047) when (flag_long='1') else '0';
	dataBufferOut(3882) <= dataBufferIn(2790) when (flag_long='1') else '0';
	dataBufferOut(3883) <= dataBufferIn(3533) when (flag_long='1') else '0';
	dataBufferOut(3884) <= dataBufferIn(4276) when (flag_long='1') else '0';
	dataBufferOut(3885) <= dataBufferIn(5019) when (flag_long='1') else '0';
	dataBufferOut(3886) <= dataBufferIn(5762) when (flag_long='1') else '0';
	dataBufferOut(3887) <= dataBufferIn( 361) when (flag_long='1') else '0';
	dataBufferOut(3888) <= dataBufferIn(1104) when (flag_long='1') else '0';
	dataBufferOut(3889) <= dataBufferIn(1847) when (flag_long='1') else '0';
	dataBufferOut(3890) <= dataBufferIn(2590) when (flag_long='1') else '0';
	dataBufferOut(3891) <= dataBufferIn(3333) when (flag_long='1') else '0';
	dataBufferOut(3892) <= dataBufferIn(4076) when (flag_long='1') else '0';
	dataBufferOut(3893) <= dataBufferIn(4819) when (flag_long='1') else '0';
	dataBufferOut(3894) <= dataBufferIn(5562) when (flag_long='1') else '0';
	dataBufferOut(3895) <= dataBufferIn( 161) when (flag_long='1') else '0';
	dataBufferOut(3896) <= dataBufferIn( 904) when (flag_long='1') else '0';
	dataBufferOut(3897) <= dataBufferIn(1647) when (flag_long='1') else '0';
	dataBufferOut(3898) <= dataBufferIn(2390) when (flag_long='1') else '0';
	dataBufferOut(3899) <= dataBufferIn(3133) when (flag_long='1') else '0';
	dataBufferOut(3900) <= dataBufferIn(3876) when (flag_long='1') else '0';
	dataBufferOut(3901) <= dataBufferIn(4619) when (flag_long='1') else '0';
	dataBufferOut(3902) <= dataBufferIn(5362) when (flag_long='1') else '0';
	dataBufferOut(3903) <= dataBufferIn(6105) when (flag_long='1') else '0';
	dataBufferOut(3904) <= dataBufferIn( 704) when (flag_long='1') else '0';
	dataBufferOut(3905) <= dataBufferIn(1447) when (flag_long='1') else '0';
	dataBufferOut(3906) <= dataBufferIn(2190) when (flag_long='1') else '0';
	dataBufferOut(3907) <= dataBufferIn(2933) when (flag_long='1') else '0';
	dataBufferOut(3908) <= dataBufferIn(3676) when (flag_long='1') else '0';
	dataBufferOut(3909) <= dataBufferIn(4419) when (flag_long='1') else '0';
	dataBufferOut(3910) <= dataBufferIn(5162) when (flag_long='1') else '0';
	dataBufferOut(3911) <= dataBufferIn(5905) when (flag_long='1') else '0';
	dataBufferOut(3912) <= dataBufferIn( 504) when (flag_long='1') else '0';
	dataBufferOut(3913) <= dataBufferIn(1247) when (flag_long='1') else '0';
	dataBufferOut(3914) <= dataBufferIn(1990) when (flag_long='1') else '0';
	dataBufferOut(3915) <= dataBufferIn(2733) when (flag_long='1') else '0';
	dataBufferOut(3916) <= dataBufferIn(3476) when (flag_long='1') else '0';
	dataBufferOut(3917) <= dataBufferIn(4219) when (flag_long='1') else '0';
	dataBufferOut(3918) <= dataBufferIn(4962) when (flag_long='1') else '0';
	dataBufferOut(3919) <= dataBufferIn(5705) when (flag_long='1') else '0';
	dataBufferOut(3920) <= dataBufferIn( 304) when (flag_long='1') else '0';
	dataBufferOut(3921) <= dataBufferIn(1047) when (flag_long='1') else '0';
	dataBufferOut(3922) <= dataBufferIn(1790) when (flag_long='1') else '0';
	dataBufferOut(3923) <= dataBufferIn(2533) when (flag_long='1') else '0';
	dataBufferOut(3924) <= dataBufferIn(3276) when (flag_long='1') else '0';
	dataBufferOut(3925) <= dataBufferIn(4019) when (flag_long='1') else '0';
	dataBufferOut(3926) <= dataBufferIn(4762) when (flag_long='1') else '0';
	dataBufferOut(3927) <= dataBufferIn(5505) when (flag_long='1') else '0';
	dataBufferOut(3928) <= dataBufferIn( 104) when (flag_long='1') else '0';
	dataBufferOut(3929) <= dataBufferIn( 847) when (flag_long='1') else '0';
	dataBufferOut(3930) <= dataBufferIn(1590) when (flag_long='1') else '0';
	dataBufferOut(3931) <= dataBufferIn(2333) when (flag_long='1') else '0';
	dataBufferOut(3932) <= dataBufferIn(3076) when (flag_long='1') else '0';
	dataBufferOut(3933) <= dataBufferIn(3819) when (flag_long='1') else '0';
	dataBufferOut(3934) <= dataBufferIn(4562) when (flag_long='1') else '0';
	dataBufferOut(3935) <= dataBufferIn(5305) when (flag_long='1') else '0';
	dataBufferOut(3936) <= dataBufferIn(6048) when (flag_long='1') else '0';
	dataBufferOut(3937) <= dataBufferIn( 647) when (flag_long='1') else '0';
	dataBufferOut(3938) <= dataBufferIn(1390) when (flag_long='1') else '0';
	dataBufferOut(3939) <= dataBufferIn(2133) when (flag_long='1') else '0';
	dataBufferOut(3940) <= dataBufferIn(2876) when (flag_long='1') else '0';
	dataBufferOut(3941) <= dataBufferIn(3619) when (flag_long='1') else '0';
	dataBufferOut(3942) <= dataBufferIn(4362) when (flag_long='1') else '0';
	dataBufferOut(3943) <= dataBufferIn(5105) when (flag_long='1') else '0';
	dataBufferOut(3944) <= dataBufferIn(5848) when (flag_long='1') else '0';
	dataBufferOut(3945) <= dataBufferIn( 447) when (flag_long='1') else '0';
	dataBufferOut(3946) <= dataBufferIn(1190) when (flag_long='1') else '0';
	dataBufferOut(3947) <= dataBufferIn(1933) when (flag_long='1') else '0';
	dataBufferOut(3948) <= dataBufferIn(2676) when (flag_long='1') else '0';
	dataBufferOut(3949) <= dataBufferIn(3419) when (flag_long='1') else '0';
	dataBufferOut(3950) <= dataBufferIn(4162) when (flag_long='1') else '0';
	dataBufferOut(3951) <= dataBufferIn(4905) when (flag_long='1') else '0';
	dataBufferOut(3952) <= dataBufferIn(5648) when (flag_long='1') else '0';
	dataBufferOut(3953) <= dataBufferIn( 247) when (flag_long='1') else '0';
	dataBufferOut(3954) <= dataBufferIn( 990) when (flag_long='1') else '0';
	dataBufferOut(3955) <= dataBufferIn(1733) when (flag_long='1') else '0';
	dataBufferOut(3956) <= dataBufferIn(2476) when (flag_long='1') else '0';
	dataBufferOut(3957) <= dataBufferIn(3219) when (flag_long='1') else '0';
	dataBufferOut(3958) <= dataBufferIn(3962) when (flag_long='1') else '0';
	dataBufferOut(3959) <= dataBufferIn(4705) when (flag_long='1') else '0';
	dataBufferOut(3960) <= dataBufferIn(5448) when (flag_long='1') else '0';
	dataBufferOut(3961) <= dataBufferIn(  47) when (flag_long='1') else '0';
	dataBufferOut(3962) <= dataBufferIn( 790) when (flag_long='1') else '0';
	dataBufferOut(3963) <= dataBufferIn(1533) when (flag_long='1') else '0';
	dataBufferOut(3964) <= dataBufferIn(2276) when (flag_long='1') else '0';
	dataBufferOut(3965) <= dataBufferIn(3019) when (flag_long='1') else '0';
	dataBufferOut(3966) <= dataBufferIn(3762) when (flag_long='1') else '0';
	dataBufferOut(3967) <= dataBufferIn(4505) when (flag_long='1') else '0';
	dataBufferOut(3968) <= dataBufferIn(5248) when (flag_long='1') else '0';
	dataBufferOut(3969) <= dataBufferIn(5991) when (flag_long='1') else '0';
	dataBufferOut(3970) <= dataBufferIn( 590) when (flag_long='1') else '0';
	dataBufferOut(3971) <= dataBufferIn(1333) when (flag_long='1') else '0';
	dataBufferOut(3972) <= dataBufferIn(2076) when (flag_long='1') else '0';
	dataBufferOut(3973) <= dataBufferIn(2819) when (flag_long='1') else '0';
	dataBufferOut(3974) <= dataBufferIn(3562) when (flag_long='1') else '0';
	dataBufferOut(3975) <= dataBufferIn(4305) when (flag_long='1') else '0';
	dataBufferOut(3976) <= dataBufferIn(5048) when (flag_long='1') else '0';
	dataBufferOut(3977) <= dataBufferIn(5791) when (flag_long='1') else '0';
	dataBufferOut(3978) <= dataBufferIn( 390) when (flag_long='1') else '0';
	dataBufferOut(3979) <= dataBufferIn(1133) when (flag_long='1') else '0';
	dataBufferOut(3980) <= dataBufferIn(1876) when (flag_long='1') else '0';
	dataBufferOut(3981) <= dataBufferIn(2619) when (flag_long='1') else '0';
	dataBufferOut(3982) <= dataBufferIn(3362) when (flag_long='1') else '0';
	dataBufferOut(3983) <= dataBufferIn(4105) when (flag_long='1') else '0';
	dataBufferOut(3984) <= dataBufferIn(4848) when (flag_long='1') else '0';
	dataBufferOut(3985) <= dataBufferIn(5591) when (flag_long='1') else '0';
	dataBufferOut(3986) <= dataBufferIn( 190) when (flag_long='1') else '0';
	dataBufferOut(3987) <= dataBufferIn( 933) when (flag_long='1') else '0';
	dataBufferOut(3988) <= dataBufferIn(1676) when (flag_long='1') else '0';
	dataBufferOut(3989) <= dataBufferIn(2419) when (flag_long='1') else '0';
	dataBufferOut(3990) <= dataBufferIn(3162) when (flag_long='1') else '0';
	dataBufferOut(3991) <= dataBufferIn(3905) when (flag_long='1') else '0';
	dataBufferOut(3992) <= dataBufferIn(4648) when (flag_long='1') else '0';
	dataBufferOut(3993) <= dataBufferIn(5391) when (flag_long='1') else '0';
	dataBufferOut(3994) <= dataBufferIn(6134) when (flag_long='1') else '0';
	dataBufferOut(3995) <= dataBufferIn( 733) when (flag_long='1') else '0';
	dataBufferOut(3996) <= dataBufferIn(1476) when (flag_long='1') else '0';
	dataBufferOut(3997) <= dataBufferIn(2219) when (flag_long='1') else '0';
	dataBufferOut(3998) <= dataBufferIn(2962) when (flag_long='1') else '0';
	dataBufferOut(3999) <= dataBufferIn(3705) when (flag_long='1') else '0';
	dataBufferOut(4000) <= dataBufferIn(4448) when (flag_long='1') else '0';
	dataBufferOut(4001) <= dataBufferIn(5191) when (flag_long='1') else '0';
	dataBufferOut(4002) <= dataBufferIn(5934) when (flag_long='1') else '0';
	dataBufferOut(4003) <= dataBufferIn( 533) when (flag_long='1') else '0';
	dataBufferOut(4004) <= dataBufferIn(1276) when (flag_long='1') else '0';
	dataBufferOut(4005) <= dataBufferIn(2019) when (flag_long='1') else '0';
	dataBufferOut(4006) <= dataBufferIn(2762) when (flag_long='1') else '0';
	dataBufferOut(4007) <= dataBufferIn(3505) when (flag_long='1') else '0';
	dataBufferOut(4008) <= dataBufferIn(4248) when (flag_long='1') else '0';
	dataBufferOut(4009) <= dataBufferIn(4991) when (flag_long='1') else '0';
	dataBufferOut(4010) <= dataBufferIn(5734) when (flag_long='1') else '0';
	dataBufferOut(4011) <= dataBufferIn( 333) when (flag_long='1') else '0';
	dataBufferOut(4012) <= dataBufferIn(1076) when (flag_long='1') else '0';
	dataBufferOut(4013) <= dataBufferIn(1819) when (flag_long='1') else '0';
	dataBufferOut(4014) <= dataBufferIn(2562) when (flag_long='1') else '0';
	dataBufferOut(4015) <= dataBufferIn(3305) when (flag_long='1') else '0';
	dataBufferOut(4016) <= dataBufferIn(4048) when (flag_long='1') else '0';
	dataBufferOut(4017) <= dataBufferIn(4791) when (flag_long='1') else '0';
	dataBufferOut(4018) <= dataBufferIn(5534) when (flag_long='1') else '0';
	dataBufferOut(4019) <= dataBufferIn( 133) when (flag_long='1') else '0';
	dataBufferOut(4020) <= dataBufferIn( 876) when (flag_long='1') else '0';
	dataBufferOut(4021) <= dataBufferIn(1619) when (flag_long='1') else '0';
	dataBufferOut(4022) <= dataBufferIn(2362) when (flag_long='1') else '0';
	dataBufferOut(4023) <= dataBufferIn(3105) when (flag_long='1') else '0';
	dataBufferOut(4024) <= dataBufferIn(3848) when (flag_long='1') else '0';
	dataBufferOut(4025) <= dataBufferIn(4591) when (flag_long='1') else '0';
	dataBufferOut(4026) <= dataBufferIn(5334) when (flag_long='1') else '0';
	dataBufferOut(4027) <= dataBufferIn(6077) when (flag_long='1') else '0';
	dataBufferOut(4028) <= dataBufferIn( 676) when (flag_long='1') else '0';
	dataBufferOut(4029) <= dataBufferIn(1419) when (flag_long='1') else '0';
	dataBufferOut(4030) <= dataBufferIn(2162) when (flag_long='1') else '0';
	dataBufferOut(4031) <= dataBufferIn(2905) when (flag_long='1') else '0';
	dataBufferOut(4032) <= dataBufferIn(3648) when (flag_long='1') else '0';
	dataBufferOut(4033) <= dataBufferIn(4391) when (flag_long='1') else '0';
	dataBufferOut(4034) <= dataBufferIn(5134) when (flag_long='1') else '0';
	dataBufferOut(4035) <= dataBufferIn(5877) when (flag_long='1') else '0';
	dataBufferOut(4036) <= dataBufferIn( 476) when (flag_long='1') else '0';
	dataBufferOut(4037) <= dataBufferIn(1219) when (flag_long='1') else '0';
	dataBufferOut(4038) <= dataBufferIn(1962) when (flag_long='1') else '0';
	dataBufferOut(4039) <= dataBufferIn(2705) when (flag_long='1') else '0';
	dataBufferOut(4040) <= dataBufferIn(3448) when (flag_long='1') else '0';
	dataBufferOut(4041) <= dataBufferIn(4191) when (flag_long='1') else '0';
	dataBufferOut(4042) <= dataBufferIn(4934) when (flag_long='1') else '0';
	dataBufferOut(4043) <= dataBufferIn(5677) when (flag_long='1') else '0';
	dataBufferOut(4044) <= dataBufferIn( 276) when (flag_long='1') else '0';
	dataBufferOut(4045) <= dataBufferIn(1019) when (flag_long='1') else '0';
	dataBufferOut(4046) <= dataBufferIn(1762) when (flag_long='1') else '0';
	dataBufferOut(4047) <= dataBufferIn(2505) when (flag_long='1') else '0';
	dataBufferOut(4048) <= dataBufferIn(3248) when (flag_long='1') else '0';
	dataBufferOut(4049) <= dataBufferIn(3991) when (flag_long='1') else '0';
	dataBufferOut(4050) <= dataBufferIn(4734) when (flag_long='1') else '0';
	dataBufferOut(4051) <= dataBufferIn(5477) when (flag_long='1') else '0';
	dataBufferOut(4052) <= dataBufferIn(  76) when (flag_long='1') else '0';
	dataBufferOut(4053) <= dataBufferIn( 819) when (flag_long='1') else '0';
	dataBufferOut(4054) <= dataBufferIn(1562) when (flag_long='1') else '0';
	dataBufferOut(4055) <= dataBufferIn(2305) when (flag_long='1') else '0';
	dataBufferOut(4056) <= dataBufferIn(3048) when (flag_long='1') else '0';
	dataBufferOut(4057) <= dataBufferIn(3791) when (flag_long='1') else '0';
	dataBufferOut(4058) <= dataBufferIn(4534) when (flag_long='1') else '0';
	dataBufferOut(4059) <= dataBufferIn(5277) when (flag_long='1') else '0';
	dataBufferOut(4060) <= dataBufferIn(6020) when (flag_long='1') else '0';
	dataBufferOut(4061) <= dataBufferIn( 619) when (flag_long='1') else '0';
	dataBufferOut(4062) <= dataBufferIn(1362) when (flag_long='1') else '0';
	dataBufferOut(4063) <= dataBufferIn(2105) when (flag_long='1') else '0';
	dataBufferOut(4064) <= dataBufferIn(2848) when (flag_long='1') else '0';
	dataBufferOut(4065) <= dataBufferIn(3591) when (flag_long='1') else '0';
	dataBufferOut(4066) <= dataBufferIn(4334) when (flag_long='1') else '0';
	dataBufferOut(4067) <= dataBufferIn(5077) when (flag_long='1') else '0';
	dataBufferOut(4068) <= dataBufferIn(5820) when (flag_long='1') else '0';
	dataBufferOut(4069) <= dataBufferIn( 419) when (flag_long='1') else '0';
	dataBufferOut(4070) <= dataBufferIn(1162) when (flag_long='1') else '0';
	dataBufferOut(4071) <= dataBufferIn(1905) when (flag_long='1') else '0';
	dataBufferOut(4072) <= dataBufferIn(2648) when (flag_long='1') else '0';
	dataBufferOut(4073) <= dataBufferIn(3391) when (flag_long='1') else '0';
	dataBufferOut(4074) <= dataBufferIn(4134) when (flag_long='1') else '0';
	dataBufferOut(4075) <= dataBufferIn(4877) when (flag_long='1') else '0';
	dataBufferOut(4076) <= dataBufferIn(5620) when (flag_long='1') else '0';
	dataBufferOut(4077) <= dataBufferIn( 219) when (flag_long='1') else '0';
	dataBufferOut(4078) <= dataBufferIn( 962) when (flag_long='1') else '0';
	dataBufferOut(4079) <= dataBufferIn(1705) when (flag_long='1') else '0';
	dataBufferOut(4080) <= dataBufferIn(2448) when (flag_long='1') else '0';
	dataBufferOut(4081) <= dataBufferIn(3191) when (flag_long='1') else '0';
	dataBufferOut(4082) <= dataBufferIn(3934) when (flag_long='1') else '0';
	dataBufferOut(4083) <= dataBufferIn(4677) when (flag_long='1') else '0';
	dataBufferOut(4084) <= dataBufferIn(5420) when (flag_long='1') else '0';
	dataBufferOut(4085) <= dataBufferIn(  19) when (flag_long='1') else '0';
	dataBufferOut(4086) <= dataBufferIn( 762) when (flag_long='1') else '0';
	dataBufferOut(4087) <= dataBufferIn(1505) when (flag_long='1') else '0';
	dataBufferOut(4088) <= dataBufferIn(2248) when (flag_long='1') else '0';
	dataBufferOut(4089) <= dataBufferIn(2991) when (flag_long='1') else '0';
	dataBufferOut(4090) <= dataBufferIn(3734) when (flag_long='1') else '0';
	dataBufferOut(4091) <= dataBufferIn(4477) when (flag_long='1') else '0';
	dataBufferOut(4092) <= dataBufferIn(5220) when (flag_long='1') else '0';
	dataBufferOut(4093) <= dataBufferIn(5963) when (flag_long='1') else '0';
	dataBufferOut(4094) <= dataBufferIn( 562) when (flag_long='1') else '0';
	dataBufferOut(4095) <= dataBufferIn(1305) when (flag_long='1') else '0';
	dataBufferOut(4096) <= dataBufferIn(2048) when (flag_long='1') else '0';
	dataBufferOut(4097) <= dataBufferIn(2791) when (flag_long='1') else '0';
	dataBufferOut(4098) <= dataBufferIn(3534) when (flag_long='1') else '0';
	dataBufferOut(4099) <= dataBufferIn(4277) when (flag_long='1') else '0';
	dataBufferOut(4100) <= dataBufferIn(5020) when (flag_long='1') else '0';
	dataBufferOut(4101) <= dataBufferIn(5763) when (flag_long='1') else '0';
	dataBufferOut(4102) <= dataBufferIn( 362) when (flag_long='1') else '0';
	dataBufferOut(4103) <= dataBufferIn(1105) when (flag_long='1') else '0';
	dataBufferOut(4104) <= dataBufferIn(1848) when (flag_long='1') else '0';
	dataBufferOut(4105) <= dataBufferIn(2591) when (flag_long='1') else '0';
	dataBufferOut(4106) <= dataBufferIn(3334) when (flag_long='1') else '0';
	dataBufferOut(4107) <= dataBufferIn(4077) when (flag_long='1') else '0';
	dataBufferOut(4108) <= dataBufferIn(4820) when (flag_long='1') else '0';
	dataBufferOut(4109) <= dataBufferIn(5563) when (flag_long='1') else '0';
	dataBufferOut(4110) <= dataBufferIn( 162) when (flag_long='1') else '0';
	dataBufferOut(4111) <= dataBufferIn( 905) when (flag_long='1') else '0';
	dataBufferOut(4112) <= dataBufferIn(1648) when (flag_long='1') else '0';
	dataBufferOut(4113) <= dataBufferIn(2391) when (flag_long='1') else '0';
	dataBufferOut(4114) <= dataBufferIn(3134) when (flag_long='1') else '0';
	dataBufferOut(4115) <= dataBufferIn(3877) when (flag_long='1') else '0';
	dataBufferOut(4116) <= dataBufferIn(4620) when (flag_long='1') else '0';
	dataBufferOut(4117) <= dataBufferIn(5363) when (flag_long='1') else '0';
	dataBufferOut(4118) <= dataBufferIn(6106) when (flag_long='1') else '0';
	dataBufferOut(4119) <= dataBufferIn( 705) when (flag_long='1') else '0';
	dataBufferOut(4120) <= dataBufferIn(1448) when (flag_long='1') else '0';
	dataBufferOut(4121) <= dataBufferIn(2191) when (flag_long='1') else '0';
	dataBufferOut(4122) <= dataBufferIn(2934) when (flag_long='1') else '0';
	dataBufferOut(4123) <= dataBufferIn(3677) when (flag_long='1') else '0';
	dataBufferOut(4124) <= dataBufferIn(4420) when (flag_long='1') else '0';
	dataBufferOut(4125) <= dataBufferIn(5163) when (flag_long='1') else '0';
	dataBufferOut(4126) <= dataBufferIn(5906) when (flag_long='1') else '0';
	dataBufferOut(4127) <= dataBufferIn( 505) when (flag_long='1') else '0';
	dataBufferOut(4128) <= dataBufferIn(1248) when (flag_long='1') else '0';
	dataBufferOut(4129) <= dataBufferIn(1991) when (flag_long='1') else '0';
	dataBufferOut(4130) <= dataBufferIn(2734) when (flag_long='1') else '0';
	dataBufferOut(4131) <= dataBufferIn(3477) when (flag_long='1') else '0';
	dataBufferOut(4132) <= dataBufferIn(4220) when (flag_long='1') else '0';
	dataBufferOut(4133) <= dataBufferIn(4963) when (flag_long='1') else '0';
	dataBufferOut(4134) <= dataBufferIn(5706) when (flag_long='1') else '0';
	dataBufferOut(4135) <= dataBufferIn( 305) when (flag_long='1') else '0';
	dataBufferOut(4136) <= dataBufferIn(1048) when (flag_long='1') else '0';
	dataBufferOut(4137) <= dataBufferIn(1791) when (flag_long='1') else '0';
	dataBufferOut(4138) <= dataBufferIn(2534) when (flag_long='1') else '0';
	dataBufferOut(4139) <= dataBufferIn(3277) when (flag_long='1') else '0';
	dataBufferOut(4140) <= dataBufferIn(4020) when (flag_long='1') else '0';
	dataBufferOut(4141) <= dataBufferIn(4763) when (flag_long='1') else '0';
	dataBufferOut(4142) <= dataBufferIn(5506) when (flag_long='1') else '0';
	dataBufferOut(4143) <= dataBufferIn( 105) when (flag_long='1') else '0';
	dataBufferOut(4144) <= dataBufferIn( 848) when (flag_long='1') else '0';
	dataBufferOut(4145) <= dataBufferIn(1591) when (flag_long='1') else '0';
	dataBufferOut(4146) <= dataBufferIn(2334) when (flag_long='1') else '0';
	dataBufferOut(4147) <= dataBufferIn(3077) when (flag_long='1') else '0';
	dataBufferOut(4148) <= dataBufferIn(3820) when (flag_long='1') else '0';
	dataBufferOut(4149) <= dataBufferIn(4563) when (flag_long='1') else '0';
	dataBufferOut(4150) <= dataBufferIn(5306) when (flag_long='1') else '0';
	dataBufferOut(4151) <= dataBufferIn(6049) when (flag_long='1') else '0';
	dataBufferOut(4152) <= dataBufferIn( 648) when (flag_long='1') else '0';
	dataBufferOut(4153) <= dataBufferIn(1391) when (flag_long='1') else '0';
	dataBufferOut(4154) <= dataBufferIn(2134) when (flag_long='1') else '0';
	dataBufferOut(4155) <= dataBufferIn(2877) when (flag_long='1') else '0';
	dataBufferOut(4156) <= dataBufferIn(3620) when (flag_long='1') else '0';
	dataBufferOut(4157) <= dataBufferIn(4363) when (flag_long='1') else '0';
	dataBufferOut(4158) <= dataBufferIn(5106) when (flag_long='1') else '0';
	dataBufferOut(4159) <= dataBufferIn(5849) when (flag_long='1') else '0';
	dataBufferOut(4160) <= dataBufferIn( 448) when (flag_long='1') else '0';
	dataBufferOut(4161) <= dataBufferIn(1191) when (flag_long='1') else '0';
	dataBufferOut(4162) <= dataBufferIn(1934) when (flag_long='1') else '0';
	dataBufferOut(4163) <= dataBufferIn(2677) when (flag_long='1') else '0';
	dataBufferOut(4164) <= dataBufferIn(3420) when (flag_long='1') else '0';
	dataBufferOut(4165) <= dataBufferIn(4163) when (flag_long='1') else '0';
	dataBufferOut(4166) <= dataBufferIn(4906) when (flag_long='1') else '0';
	dataBufferOut(4167) <= dataBufferIn(5649) when (flag_long='1') else '0';
	dataBufferOut(4168) <= dataBufferIn( 248) when (flag_long='1') else '0';
	dataBufferOut(4169) <= dataBufferIn( 991) when (flag_long='1') else '0';
	dataBufferOut(4170) <= dataBufferIn(1734) when (flag_long='1') else '0';
	dataBufferOut(4171) <= dataBufferIn(2477) when (flag_long='1') else '0';
	dataBufferOut(4172) <= dataBufferIn(3220) when (flag_long='1') else '0';
	dataBufferOut(4173) <= dataBufferIn(3963) when (flag_long='1') else '0';
	dataBufferOut(4174) <= dataBufferIn(4706) when (flag_long='1') else '0';
	dataBufferOut(4175) <= dataBufferIn(5449) when (flag_long='1') else '0';
	dataBufferOut(4176) <= dataBufferIn(  48) when (flag_long='1') else '0';
	dataBufferOut(4177) <= dataBufferIn( 791) when (flag_long='1') else '0';
	dataBufferOut(4178) <= dataBufferIn(1534) when (flag_long='1') else '0';
	dataBufferOut(4179) <= dataBufferIn(2277) when (flag_long='1') else '0';
	dataBufferOut(4180) <= dataBufferIn(3020) when (flag_long='1') else '0';
	dataBufferOut(4181) <= dataBufferIn(3763) when (flag_long='1') else '0';
	dataBufferOut(4182) <= dataBufferIn(4506) when (flag_long='1') else '0';
	dataBufferOut(4183) <= dataBufferIn(5249) when (flag_long='1') else '0';
	dataBufferOut(4184) <= dataBufferIn(5992) when (flag_long='1') else '0';
	dataBufferOut(4185) <= dataBufferIn( 591) when (flag_long='1') else '0';
	dataBufferOut(4186) <= dataBufferIn(1334) when (flag_long='1') else '0';
	dataBufferOut(4187) <= dataBufferIn(2077) when (flag_long='1') else '0';
	dataBufferOut(4188) <= dataBufferIn(2820) when (flag_long='1') else '0';
	dataBufferOut(4189) <= dataBufferIn(3563) when (flag_long='1') else '0';
	dataBufferOut(4190) <= dataBufferIn(4306) when (flag_long='1') else '0';
	dataBufferOut(4191) <= dataBufferIn(5049) when (flag_long='1') else '0';
	dataBufferOut(4192) <= dataBufferIn(5792) when (flag_long='1') else '0';
	dataBufferOut(4193) <= dataBufferIn( 391) when (flag_long='1') else '0';
	dataBufferOut(4194) <= dataBufferIn(1134) when (flag_long='1') else '0';
	dataBufferOut(4195) <= dataBufferIn(1877) when (flag_long='1') else '0';
	dataBufferOut(4196) <= dataBufferIn(2620) when (flag_long='1') else '0';
	dataBufferOut(4197) <= dataBufferIn(3363) when (flag_long='1') else '0';
	dataBufferOut(4198) <= dataBufferIn(4106) when (flag_long='1') else '0';
	dataBufferOut(4199) <= dataBufferIn(4849) when (flag_long='1') else '0';
	dataBufferOut(4200) <= dataBufferIn(5592) when (flag_long='1') else '0';
	dataBufferOut(4201) <= dataBufferIn( 191) when (flag_long='1') else '0';
	dataBufferOut(4202) <= dataBufferIn( 934) when (flag_long='1') else '0';
	dataBufferOut(4203) <= dataBufferIn(1677) when (flag_long='1') else '0';
	dataBufferOut(4204) <= dataBufferIn(2420) when (flag_long='1') else '0';
	dataBufferOut(4205) <= dataBufferIn(3163) when (flag_long='1') else '0';
	dataBufferOut(4206) <= dataBufferIn(3906) when (flag_long='1') else '0';
	dataBufferOut(4207) <= dataBufferIn(4649) when (flag_long='1') else '0';
	dataBufferOut(4208) <= dataBufferIn(5392) when (flag_long='1') else '0';
	dataBufferOut(4209) <= dataBufferIn(6135) when (flag_long='1') else '0';
	dataBufferOut(4210) <= dataBufferIn( 734) when (flag_long='1') else '0';
	dataBufferOut(4211) <= dataBufferIn(1477) when (flag_long='1') else '0';
	dataBufferOut(4212) <= dataBufferIn(2220) when (flag_long='1') else '0';
	dataBufferOut(4213) <= dataBufferIn(2963) when (flag_long='1') else '0';
	dataBufferOut(4214) <= dataBufferIn(3706) when (flag_long='1') else '0';
	dataBufferOut(4215) <= dataBufferIn(4449) when (flag_long='1') else '0';
	dataBufferOut(4216) <= dataBufferIn(5192) when (flag_long='1') else '0';
	dataBufferOut(4217) <= dataBufferIn(5935) when (flag_long='1') else '0';
	dataBufferOut(4218) <= dataBufferIn( 534) when (flag_long='1') else '0';
	dataBufferOut(4219) <= dataBufferIn(1277) when (flag_long='1') else '0';
	dataBufferOut(4220) <= dataBufferIn(2020) when (flag_long='1') else '0';
	dataBufferOut(4221) <= dataBufferIn(2763) when (flag_long='1') else '0';
	dataBufferOut(4222) <= dataBufferIn(3506) when (flag_long='1') else '0';
	dataBufferOut(4223) <= dataBufferIn(4249) when (flag_long='1') else '0';
	dataBufferOut(4224) <= dataBufferIn(4992) when (flag_long='1') else '0';
	dataBufferOut(4225) <= dataBufferIn(5735) when (flag_long='1') else '0';
	dataBufferOut(4226) <= dataBufferIn( 334) when (flag_long='1') else '0';
	dataBufferOut(4227) <= dataBufferIn(1077) when (flag_long='1') else '0';
	dataBufferOut(4228) <= dataBufferIn(1820) when (flag_long='1') else '0';
	dataBufferOut(4229) <= dataBufferIn(2563) when (flag_long='1') else '0';
	dataBufferOut(4230) <= dataBufferIn(3306) when (flag_long='1') else '0';
	dataBufferOut(4231) <= dataBufferIn(4049) when (flag_long='1') else '0';
	dataBufferOut(4232) <= dataBufferIn(4792) when (flag_long='1') else '0';
	dataBufferOut(4233) <= dataBufferIn(5535) when (flag_long='1') else '0';
	dataBufferOut(4234) <= dataBufferIn( 134) when (flag_long='1') else '0';
	dataBufferOut(4235) <= dataBufferIn( 877) when (flag_long='1') else '0';
	dataBufferOut(4236) <= dataBufferIn(1620) when (flag_long='1') else '0';
	dataBufferOut(4237) <= dataBufferIn(2363) when (flag_long='1') else '0';
	dataBufferOut(4238) <= dataBufferIn(3106) when (flag_long='1') else '0';
	dataBufferOut(4239) <= dataBufferIn(3849) when (flag_long='1') else '0';
	dataBufferOut(4240) <= dataBufferIn(4592) when (flag_long='1') else '0';
	dataBufferOut(4241) <= dataBufferIn(5335) when (flag_long='1') else '0';
	dataBufferOut(4242) <= dataBufferIn(6078) when (flag_long='1') else '0';
	dataBufferOut(4243) <= dataBufferIn( 677) when (flag_long='1') else '0';
	dataBufferOut(4244) <= dataBufferIn(1420) when (flag_long='1') else '0';
	dataBufferOut(4245) <= dataBufferIn(2163) when (flag_long='1') else '0';
	dataBufferOut(4246) <= dataBufferIn(2906) when (flag_long='1') else '0';
	dataBufferOut(4247) <= dataBufferIn(3649) when (flag_long='1') else '0';
	dataBufferOut(4248) <= dataBufferIn(4392) when (flag_long='1') else '0';
	dataBufferOut(4249) <= dataBufferIn(5135) when (flag_long='1') else '0';
	dataBufferOut(4250) <= dataBufferIn(5878) when (flag_long='1') else '0';
	dataBufferOut(4251) <= dataBufferIn( 477) when (flag_long='1') else '0';
	dataBufferOut(4252) <= dataBufferIn(1220) when (flag_long='1') else '0';
	dataBufferOut(4253) <= dataBufferIn(1963) when (flag_long='1') else '0';
	dataBufferOut(4254) <= dataBufferIn(2706) when (flag_long='1') else '0';
	dataBufferOut(4255) <= dataBufferIn(3449) when (flag_long='1') else '0';
	dataBufferOut(4256) <= dataBufferIn(4192) when (flag_long='1') else '0';
	dataBufferOut(4257) <= dataBufferIn(4935) when (flag_long='1') else '0';
	dataBufferOut(4258) <= dataBufferIn(5678) when (flag_long='1') else '0';
	dataBufferOut(4259) <= dataBufferIn( 277) when (flag_long='1') else '0';
	dataBufferOut(4260) <= dataBufferIn(1020) when (flag_long='1') else '0';
	dataBufferOut(4261) <= dataBufferIn(1763) when (flag_long='1') else '0';
	dataBufferOut(4262) <= dataBufferIn(2506) when (flag_long='1') else '0';
	dataBufferOut(4263) <= dataBufferIn(3249) when (flag_long='1') else '0';
	dataBufferOut(4264) <= dataBufferIn(3992) when (flag_long='1') else '0';
	dataBufferOut(4265) <= dataBufferIn(4735) when (flag_long='1') else '0';
	dataBufferOut(4266) <= dataBufferIn(5478) when (flag_long='1') else '0';
	dataBufferOut(4267) <= dataBufferIn(  77) when (flag_long='1') else '0';
	dataBufferOut(4268) <= dataBufferIn( 820) when (flag_long='1') else '0';
	dataBufferOut(4269) <= dataBufferIn(1563) when (flag_long='1') else '0';
	dataBufferOut(4270) <= dataBufferIn(2306) when (flag_long='1') else '0';
	dataBufferOut(4271) <= dataBufferIn(3049) when (flag_long='1') else '0';
	dataBufferOut(4272) <= dataBufferIn(3792) when (flag_long='1') else '0';
	dataBufferOut(4273) <= dataBufferIn(4535) when (flag_long='1') else '0';
	dataBufferOut(4274) <= dataBufferIn(5278) when (flag_long='1') else '0';
	dataBufferOut(4275) <= dataBufferIn(6021) when (flag_long='1') else '0';
	dataBufferOut(4276) <= dataBufferIn( 620) when (flag_long='1') else '0';
	dataBufferOut(4277) <= dataBufferIn(1363) when (flag_long='1') else '0';
	dataBufferOut(4278) <= dataBufferIn(2106) when (flag_long='1') else '0';
	dataBufferOut(4279) <= dataBufferIn(2849) when (flag_long='1') else '0';
	dataBufferOut(4280) <= dataBufferIn(3592) when (flag_long='1') else '0';
	dataBufferOut(4281) <= dataBufferIn(4335) when (flag_long='1') else '0';
	dataBufferOut(4282) <= dataBufferIn(5078) when (flag_long='1') else '0';
	dataBufferOut(4283) <= dataBufferIn(5821) when (flag_long='1') else '0';
	dataBufferOut(4284) <= dataBufferIn( 420) when (flag_long='1') else '0';
	dataBufferOut(4285) <= dataBufferIn(1163) when (flag_long='1') else '0';
	dataBufferOut(4286) <= dataBufferIn(1906) when (flag_long='1') else '0';
	dataBufferOut(4287) <= dataBufferIn(2649) when (flag_long='1') else '0';
	dataBufferOut(4288) <= dataBufferIn(3392) when (flag_long='1') else '0';
	dataBufferOut(4289) <= dataBufferIn(4135) when (flag_long='1') else '0';
	dataBufferOut(4290) <= dataBufferIn(4878) when (flag_long='1') else '0';
	dataBufferOut(4291) <= dataBufferIn(5621) when (flag_long='1') else '0';
	dataBufferOut(4292) <= dataBufferIn( 220) when (flag_long='1') else '0';
	dataBufferOut(4293) <= dataBufferIn( 963) when (flag_long='1') else '0';
	dataBufferOut(4294) <= dataBufferIn(1706) when (flag_long='1') else '0';
	dataBufferOut(4295) <= dataBufferIn(2449) when (flag_long='1') else '0';
	dataBufferOut(4296) <= dataBufferIn(3192) when (flag_long='1') else '0';
	dataBufferOut(4297) <= dataBufferIn(3935) when (flag_long='1') else '0';
	dataBufferOut(4298) <= dataBufferIn(4678) when (flag_long='1') else '0';
	dataBufferOut(4299) <= dataBufferIn(5421) when (flag_long='1') else '0';
	dataBufferOut(4300) <= dataBufferIn(  20) when (flag_long='1') else '0';
	dataBufferOut(4301) <= dataBufferIn( 763) when (flag_long='1') else '0';
	dataBufferOut(4302) <= dataBufferIn(1506) when (flag_long='1') else '0';
	dataBufferOut(4303) <= dataBufferIn(2249) when (flag_long='1') else '0';
	dataBufferOut(4304) <= dataBufferIn(2992) when (flag_long='1') else '0';
	dataBufferOut(4305) <= dataBufferIn(3735) when (flag_long='1') else '0';
	dataBufferOut(4306) <= dataBufferIn(4478) when (flag_long='1') else '0';
	dataBufferOut(4307) <= dataBufferIn(5221) when (flag_long='1') else '0';
	dataBufferOut(4308) <= dataBufferIn(5964) when (flag_long='1') else '0';
	dataBufferOut(4309) <= dataBufferIn( 563) when (flag_long='1') else '0';
	dataBufferOut(4310) <= dataBufferIn(1306) when (flag_long='1') else '0';
	dataBufferOut(4311) <= dataBufferIn(2049) when (flag_long='1') else '0';
	dataBufferOut(4312) <= dataBufferIn(2792) when (flag_long='1') else '0';
	dataBufferOut(4313) <= dataBufferIn(3535) when (flag_long='1') else '0';
	dataBufferOut(4314) <= dataBufferIn(4278) when (flag_long='1') else '0';
	dataBufferOut(4315) <= dataBufferIn(5021) when (flag_long='1') else '0';
	dataBufferOut(4316) <= dataBufferIn(5764) when (flag_long='1') else '0';
	dataBufferOut(4317) <= dataBufferIn( 363) when (flag_long='1') else '0';
	dataBufferOut(4318) <= dataBufferIn(1106) when (flag_long='1') else '0';
	dataBufferOut(4319) <= dataBufferIn(1849) when (flag_long='1') else '0';
	dataBufferOut(4320) <= dataBufferIn(2592) when (flag_long='1') else '0';
	dataBufferOut(4321) <= dataBufferIn(3335) when (flag_long='1') else '0';
	dataBufferOut(4322) <= dataBufferIn(4078) when (flag_long='1') else '0';
	dataBufferOut(4323) <= dataBufferIn(4821) when (flag_long='1') else '0';
	dataBufferOut(4324) <= dataBufferIn(5564) when (flag_long='1') else '0';
	dataBufferOut(4325) <= dataBufferIn( 163) when (flag_long='1') else '0';
	dataBufferOut(4326) <= dataBufferIn( 906) when (flag_long='1') else '0';
	dataBufferOut(4327) <= dataBufferIn(1649) when (flag_long='1') else '0';
	dataBufferOut(4328) <= dataBufferIn(2392) when (flag_long='1') else '0';
	dataBufferOut(4329) <= dataBufferIn(3135) when (flag_long='1') else '0';
	dataBufferOut(4330) <= dataBufferIn(3878) when (flag_long='1') else '0';
	dataBufferOut(4331) <= dataBufferIn(4621) when (flag_long='1') else '0';
	dataBufferOut(4332) <= dataBufferIn(5364) when (flag_long='1') else '0';
	dataBufferOut(4333) <= dataBufferIn(6107) when (flag_long='1') else '0';
	dataBufferOut(4334) <= dataBufferIn( 706) when (flag_long='1') else '0';
	dataBufferOut(4335) <= dataBufferIn(1449) when (flag_long='1') else '0';
	dataBufferOut(4336) <= dataBufferIn(2192) when (flag_long='1') else '0';
	dataBufferOut(4337) <= dataBufferIn(2935) when (flag_long='1') else '0';
	dataBufferOut(4338) <= dataBufferIn(3678) when (flag_long='1') else '0';
	dataBufferOut(4339) <= dataBufferIn(4421) when (flag_long='1') else '0';
	dataBufferOut(4340) <= dataBufferIn(5164) when (flag_long='1') else '0';
	dataBufferOut(4341) <= dataBufferIn(5907) when (flag_long='1') else '0';
	dataBufferOut(4342) <= dataBufferIn( 506) when (flag_long='1') else '0';
	dataBufferOut(4343) <= dataBufferIn(1249) when (flag_long='1') else '0';
	dataBufferOut(4344) <= dataBufferIn(1992) when (flag_long='1') else '0';
	dataBufferOut(4345) <= dataBufferIn(2735) when (flag_long='1') else '0';
	dataBufferOut(4346) <= dataBufferIn(3478) when (flag_long='1') else '0';
	dataBufferOut(4347) <= dataBufferIn(4221) when (flag_long='1') else '0';
	dataBufferOut(4348) <= dataBufferIn(4964) when (flag_long='1') else '0';
	dataBufferOut(4349) <= dataBufferIn(5707) when (flag_long='1') else '0';
	dataBufferOut(4350) <= dataBufferIn( 306) when (flag_long='1') else '0';
	dataBufferOut(4351) <= dataBufferIn(1049) when (flag_long='1') else '0';
	dataBufferOut(4352) <= dataBufferIn(1792) when (flag_long='1') else '0';
	dataBufferOut(4353) <= dataBufferIn(2535) when (flag_long='1') else '0';
	dataBufferOut(4354) <= dataBufferIn(3278) when (flag_long='1') else '0';
	dataBufferOut(4355) <= dataBufferIn(4021) when (flag_long='1') else '0';
	dataBufferOut(4356) <= dataBufferIn(4764) when (flag_long='1') else '0';
	dataBufferOut(4357) <= dataBufferIn(5507) when (flag_long='1') else '0';
	dataBufferOut(4358) <= dataBufferIn( 106) when (flag_long='1') else '0';
	dataBufferOut(4359) <= dataBufferIn( 849) when (flag_long='1') else '0';
	dataBufferOut(4360) <= dataBufferIn(1592) when (flag_long='1') else '0';
	dataBufferOut(4361) <= dataBufferIn(2335) when (flag_long='1') else '0';
	dataBufferOut(4362) <= dataBufferIn(3078) when (flag_long='1') else '0';
	dataBufferOut(4363) <= dataBufferIn(3821) when (flag_long='1') else '0';
	dataBufferOut(4364) <= dataBufferIn(4564) when (flag_long='1') else '0';
	dataBufferOut(4365) <= dataBufferIn(5307) when (flag_long='1') else '0';
	dataBufferOut(4366) <= dataBufferIn(6050) when (flag_long='1') else '0';
	dataBufferOut(4367) <= dataBufferIn( 649) when (flag_long='1') else '0';
	dataBufferOut(4368) <= dataBufferIn(1392) when (flag_long='1') else '0';
	dataBufferOut(4369) <= dataBufferIn(2135) when (flag_long='1') else '0';
	dataBufferOut(4370) <= dataBufferIn(2878) when (flag_long='1') else '0';
	dataBufferOut(4371) <= dataBufferIn(3621) when (flag_long='1') else '0';
	dataBufferOut(4372) <= dataBufferIn(4364) when (flag_long='1') else '0';
	dataBufferOut(4373) <= dataBufferIn(5107) when (flag_long='1') else '0';
	dataBufferOut(4374) <= dataBufferIn(5850) when (flag_long='1') else '0';
	dataBufferOut(4375) <= dataBufferIn( 449) when (flag_long='1') else '0';
	dataBufferOut(4376) <= dataBufferIn(1192) when (flag_long='1') else '0';
	dataBufferOut(4377) <= dataBufferIn(1935) when (flag_long='1') else '0';
	dataBufferOut(4378) <= dataBufferIn(2678) when (flag_long='1') else '0';
	dataBufferOut(4379) <= dataBufferIn(3421) when (flag_long='1') else '0';
	dataBufferOut(4380) <= dataBufferIn(4164) when (flag_long='1') else '0';
	dataBufferOut(4381) <= dataBufferIn(4907) when (flag_long='1') else '0';
	dataBufferOut(4382) <= dataBufferIn(5650) when (flag_long='1') else '0';
	dataBufferOut(4383) <= dataBufferIn( 249) when (flag_long='1') else '0';
	dataBufferOut(4384) <= dataBufferIn( 992) when (flag_long='1') else '0';
	dataBufferOut(4385) <= dataBufferIn(1735) when (flag_long='1') else '0';
	dataBufferOut(4386) <= dataBufferIn(2478) when (flag_long='1') else '0';
	dataBufferOut(4387) <= dataBufferIn(3221) when (flag_long='1') else '0';
	dataBufferOut(4388) <= dataBufferIn(3964) when (flag_long='1') else '0';
	dataBufferOut(4389) <= dataBufferIn(4707) when (flag_long='1') else '0';
	dataBufferOut(4390) <= dataBufferIn(5450) when (flag_long='1') else '0';
	dataBufferOut(4391) <= dataBufferIn(  49) when (flag_long='1') else '0';
	dataBufferOut(4392) <= dataBufferIn( 792) when (flag_long='1') else '0';
	dataBufferOut(4393) <= dataBufferIn(1535) when (flag_long='1') else '0';
	dataBufferOut(4394) <= dataBufferIn(2278) when (flag_long='1') else '0';
	dataBufferOut(4395) <= dataBufferIn(3021) when (flag_long='1') else '0';
	dataBufferOut(4396) <= dataBufferIn(3764) when (flag_long='1') else '0';
	dataBufferOut(4397) <= dataBufferIn(4507) when (flag_long='1') else '0';
	dataBufferOut(4398) <= dataBufferIn(5250) when (flag_long='1') else '0';
	dataBufferOut(4399) <= dataBufferIn(5993) when (flag_long='1') else '0';
	dataBufferOut(4400) <= dataBufferIn( 592) when (flag_long='1') else '0';
	dataBufferOut(4401) <= dataBufferIn(1335) when (flag_long='1') else '0';
	dataBufferOut(4402) <= dataBufferIn(2078) when (flag_long='1') else '0';
	dataBufferOut(4403) <= dataBufferIn(2821) when (flag_long='1') else '0';
	dataBufferOut(4404) <= dataBufferIn(3564) when (flag_long='1') else '0';
	dataBufferOut(4405) <= dataBufferIn(4307) when (flag_long='1') else '0';
	dataBufferOut(4406) <= dataBufferIn(5050) when (flag_long='1') else '0';
	dataBufferOut(4407) <= dataBufferIn(5793) when (flag_long='1') else '0';
	dataBufferOut(4408) <= dataBufferIn( 392) when (flag_long='1') else '0';
	dataBufferOut(4409) <= dataBufferIn(1135) when (flag_long='1') else '0';
	dataBufferOut(4410) <= dataBufferIn(1878) when (flag_long='1') else '0';
	dataBufferOut(4411) <= dataBufferIn(2621) when (flag_long='1') else '0';
	dataBufferOut(4412) <= dataBufferIn(3364) when (flag_long='1') else '0';
	dataBufferOut(4413) <= dataBufferIn(4107) when (flag_long='1') else '0';
	dataBufferOut(4414) <= dataBufferIn(4850) when (flag_long='1') else '0';
	dataBufferOut(4415) <= dataBufferIn(5593) when (flag_long='1') else '0';
	dataBufferOut(4416) <= dataBufferIn( 192) when (flag_long='1') else '0';
	dataBufferOut(4417) <= dataBufferIn( 935) when (flag_long='1') else '0';
	dataBufferOut(4418) <= dataBufferIn(1678) when (flag_long='1') else '0';
	dataBufferOut(4419) <= dataBufferIn(2421) when (flag_long='1') else '0';
	dataBufferOut(4420) <= dataBufferIn(3164) when (flag_long='1') else '0';
	dataBufferOut(4421) <= dataBufferIn(3907) when (flag_long='1') else '0';
	dataBufferOut(4422) <= dataBufferIn(4650) when (flag_long='1') else '0';
	dataBufferOut(4423) <= dataBufferIn(5393) when (flag_long='1') else '0';
	dataBufferOut(4424) <= dataBufferIn(6136) when (flag_long='1') else '0';
	dataBufferOut(4425) <= dataBufferIn( 735) when (flag_long='1') else '0';
	dataBufferOut(4426) <= dataBufferIn(1478) when (flag_long='1') else '0';
	dataBufferOut(4427) <= dataBufferIn(2221) when (flag_long='1') else '0';
	dataBufferOut(4428) <= dataBufferIn(2964) when (flag_long='1') else '0';
	dataBufferOut(4429) <= dataBufferIn(3707) when (flag_long='1') else '0';
	dataBufferOut(4430) <= dataBufferIn(4450) when (flag_long='1') else '0';
	dataBufferOut(4431) <= dataBufferIn(5193) when (flag_long='1') else '0';
	dataBufferOut(4432) <= dataBufferIn(5936) when (flag_long='1') else '0';
	dataBufferOut(4433) <= dataBufferIn( 535) when (flag_long='1') else '0';
	dataBufferOut(4434) <= dataBufferIn(1278) when (flag_long='1') else '0';
	dataBufferOut(4435) <= dataBufferIn(2021) when (flag_long='1') else '0';
	dataBufferOut(4436) <= dataBufferIn(2764) when (flag_long='1') else '0';
	dataBufferOut(4437) <= dataBufferIn(3507) when (flag_long='1') else '0';
	dataBufferOut(4438) <= dataBufferIn(4250) when (flag_long='1') else '0';
	dataBufferOut(4439) <= dataBufferIn(4993) when (flag_long='1') else '0';
	dataBufferOut(4440) <= dataBufferIn(5736) when (flag_long='1') else '0';
	dataBufferOut(4441) <= dataBufferIn( 335) when (flag_long='1') else '0';
	dataBufferOut(4442) <= dataBufferIn(1078) when (flag_long='1') else '0';
	dataBufferOut(4443) <= dataBufferIn(1821) when (flag_long='1') else '0';
	dataBufferOut(4444) <= dataBufferIn(2564) when (flag_long='1') else '0';
	dataBufferOut(4445) <= dataBufferIn(3307) when (flag_long='1') else '0';
	dataBufferOut(4446) <= dataBufferIn(4050) when (flag_long='1') else '0';
	dataBufferOut(4447) <= dataBufferIn(4793) when (flag_long='1') else '0';
	dataBufferOut(4448) <= dataBufferIn(5536) when (flag_long='1') else '0';
	dataBufferOut(4449) <= dataBufferIn( 135) when (flag_long='1') else '0';
	dataBufferOut(4450) <= dataBufferIn( 878) when (flag_long='1') else '0';
	dataBufferOut(4451) <= dataBufferIn(1621) when (flag_long='1') else '0';
	dataBufferOut(4452) <= dataBufferIn(2364) when (flag_long='1') else '0';
	dataBufferOut(4453) <= dataBufferIn(3107) when (flag_long='1') else '0';
	dataBufferOut(4454) <= dataBufferIn(3850) when (flag_long='1') else '0';
	dataBufferOut(4455) <= dataBufferIn(4593) when (flag_long='1') else '0';
	dataBufferOut(4456) <= dataBufferIn(5336) when (flag_long='1') else '0';
	dataBufferOut(4457) <= dataBufferIn(6079) when (flag_long='1') else '0';
	dataBufferOut(4458) <= dataBufferIn( 678) when (flag_long='1') else '0';
	dataBufferOut(4459) <= dataBufferIn(1421) when (flag_long='1') else '0';
	dataBufferOut(4460) <= dataBufferIn(2164) when (flag_long='1') else '0';
	dataBufferOut(4461) <= dataBufferIn(2907) when (flag_long='1') else '0';
	dataBufferOut(4462) <= dataBufferIn(3650) when (flag_long='1') else '0';
	dataBufferOut(4463) <= dataBufferIn(4393) when (flag_long='1') else '0';
	dataBufferOut(4464) <= dataBufferIn(5136) when (flag_long='1') else '0';
	dataBufferOut(4465) <= dataBufferIn(5879) when (flag_long='1') else '0';
	dataBufferOut(4466) <= dataBufferIn( 478) when (flag_long='1') else '0';
	dataBufferOut(4467) <= dataBufferIn(1221) when (flag_long='1') else '0';
	dataBufferOut(4468) <= dataBufferIn(1964) when (flag_long='1') else '0';
	dataBufferOut(4469) <= dataBufferIn(2707) when (flag_long='1') else '0';
	dataBufferOut(4470) <= dataBufferIn(3450) when (flag_long='1') else '0';
	dataBufferOut(4471) <= dataBufferIn(4193) when (flag_long='1') else '0';
	dataBufferOut(4472) <= dataBufferIn(4936) when (flag_long='1') else '0';
	dataBufferOut(4473) <= dataBufferIn(5679) when (flag_long='1') else '0';
	dataBufferOut(4474) <= dataBufferIn( 278) when (flag_long='1') else '0';
	dataBufferOut(4475) <= dataBufferIn(1021) when (flag_long='1') else '0';
	dataBufferOut(4476) <= dataBufferIn(1764) when (flag_long='1') else '0';
	dataBufferOut(4477) <= dataBufferIn(2507) when (flag_long='1') else '0';
	dataBufferOut(4478) <= dataBufferIn(3250) when (flag_long='1') else '0';
	dataBufferOut(4479) <= dataBufferIn(3993) when (flag_long='1') else '0';
	dataBufferOut(4480) <= dataBufferIn(4736) when (flag_long='1') else '0';
	dataBufferOut(4481) <= dataBufferIn(5479) when (flag_long='1') else '0';
	dataBufferOut(4482) <= dataBufferIn(  78) when (flag_long='1') else '0';
	dataBufferOut(4483) <= dataBufferIn( 821) when (flag_long='1') else '0';
	dataBufferOut(4484) <= dataBufferIn(1564) when (flag_long='1') else '0';
	dataBufferOut(4485) <= dataBufferIn(2307) when (flag_long='1') else '0';
	dataBufferOut(4486) <= dataBufferIn(3050) when (flag_long='1') else '0';
	dataBufferOut(4487) <= dataBufferIn(3793) when (flag_long='1') else '0';
	dataBufferOut(4488) <= dataBufferIn(4536) when (flag_long='1') else '0';
	dataBufferOut(4489) <= dataBufferIn(5279) when (flag_long='1') else '0';
	dataBufferOut(4490) <= dataBufferIn(6022) when (flag_long='1') else '0';
	dataBufferOut(4491) <= dataBufferIn( 621) when (flag_long='1') else '0';
	dataBufferOut(4492) <= dataBufferIn(1364) when (flag_long='1') else '0';
	dataBufferOut(4493) <= dataBufferIn(2107) when (flag_long='1') else '0';
	dataBufferOut(4494) <= dataBufferIn(2850) when (flag_long='1') else '0';
	dataBufferOut(4495) <= dataBufferIn(3593) when (flag_long='1') else '0';
	dataBufferOut(4496) <= dataBufferIn(4336) when (flag_long='1') else '0';
	dataBufferOut(4497) <= dataBufferIn(5079) when (flag_long='1') else '0';
	dataBufferOut(4498) <= dataBufferIn(5822) when (flag_long='1') else '0';
	dataBufferOut(4499) <= dataBufferIn( 421) when (flag_long='1') else '0';
	dataBufferOut(4500) <= dataBufferIn(1164) when (flag_long='1') else '0';
	dataBufferOut(4501) <= dataBufferIn(1907) when (flag_long='1') else '0';
	dataBufferOut(4502) <= dataBufferIn(2650) when (flag_long='1') else '0';
	dataBufferOut(4503) <= dataBufferIn(3393) when (flag_long='1') else '0';
	dataBufferOut(4504) <= dataBufferIn(4136) when (flag_long='1') else '0';
	dataBufferOut(4505) <= dataBufferIn(4879) when (flag_long='1') else '0';
	dataBufferOut(4506) <= dataBufferIn(5622) when (flag_long='1') else '0';
	dataBufferOut(4507) <= dataBufferIn( 221) when (flag_long='1') else '0';
	dataBufferOut(4508) <= dataBufferIn( 964) when (flag_long='1') else '0';
	dataBufferOut(4509) <= dataBufferIn(1707) when (flag_long='1') else '0';
	dataBufferOut(4510) <= dataBufferIn(2450) when (flag_long='1') else '0';
	dataBufferOut(4511) <= dataBufferIn(3193) when (flag_long='1') else '0';
	dataBufferOut(4512) <= dataBufferIn(3936) when (flag_long='1') else '0';
	dataBufferOut(4513) <= dataBufferIn(4679) when (flag_long='1') else '0';
	dataBufferOut(4514) <= dataBufferIn(5422) when (flag_long='1') else '0';
	dataBufferOut(4515) <= dataBufferIn(  21) when (flag_long='1') else '0';
	dataBufferOut(4516) <= dataBufferIn( 764) when (flag_long='1') else '0';
	dataBufferOut(4517) <= dataBufferIn(1507) when (flag_long='1') else '0';
	dataBufferOut(4518) <= dataBufferIn(2250) when (flag_long='1') else '0';
	dataBufferOut(4519) <= dataBufferIn(2993) when (flag_long='1') else '0';
	dataBufferOut(4520) <= dataBufferIn(3736) when (flag_long='1') else '0';
	dataBufferOut(4521) <= dataBufferIn(4479) when (flag_long='1') else '0';
	dataBufferOut(4522) <= dataBufferIn(5222) when (flag_long='1') else '0';
	dataBufferOut(4523) <= dataBufferIn(5965) when (flag_long='1') else '0';
	dataBufferOut(4524) <= dataBufferIn( 564) when (flag_long='1') else '0';
	dataBufferOut(4525) <= dataBufferIn(1307) when (flag_long='1') else '0';
	dataBufferOut(4526) <= dataBufferIn(2050) when (flag_long='1') else '0';
	dataBufferOut(4527) <= dataBufferIn(2793) when (flag_long='1') else '0';
	dataBufferOut(4528) <= dataBufferIn(3536) when (flag_long='1') else '0';
	dataBufferOut(4529) <= dataBufferIn(4279) when (flag_long='1') else '0';
	dataBufferOut(4530) <= dataBufferIn(5022) when (flag_long='1') else '0';
	dataBufferOut(4531) <= dataBufferIn(5765) when (flag_long='1') else '0';
	dataBufferOut(4532) <= dataBufferIn( 364) when (flag_long='1') else '0';
	dataBufferOut(4533) <= dataBufferIn(1107) when (flag_long='1') else '0';
	dataBufferOut(4534) <= dataBufferIn(1850) when (flag_long='1') else '0';
	dataBufferOut(4535) <= dataBufferIn(2593) when (flag_long='1') else '0';
	dataBufferOut(4536) <= dataBufferIn(3336) when (flag_long='1') else '0';
	dataBufferOut(4537) <= dataBufferIn(4079) when (flag_long='1') else '0';
	dataBufferOut(4538) <= dataBufferIn(4822) when (flag_long='1') else '0';
	dataBufferOut(4539) <= dataBufferIn(5565) when (flag_long='1') else '0';
	dataBufferOut(4540) <= dataBufferIn( 164) when (flag_long='1') else '0';
	dataBufferOut(4541) <= dataBufferIn( 907) when (flag_long='1') else '0';
	dataBufferOut(4542) <= dataBufferIn(1650) when (flag_long='1') else '0';
	dataBufferOut(4543) <= dataBufferIn(2393) when (flag_long='1') else '0';
	dataBufferOut(4544) <= dataBufferIn(3136) when (flag_long='1') else '0';
	dataBufferOut(4545) <= dataBufferIn(3879) when (flag_long='1') else '0';
	dataBufferOut(4546) <= dataBufferIn(4622) when (flag_long='1') else '0';
	dataBufferOut(4547) <= dataBufferIn(5365) when (flag_long='1') else '0';
	dataBufferOut(4548) <= dataBufferIn(6108) when (flag_long='1') else '0';
	dataBufferOut(4549) <= dataBufferIn( 707) when (flag_long='1') else '0';
	dataBufferOut(4550) <= dataBufferIn(1450) when (flag_long='1') else '0';
	dataBufferOut(4551) <= dataBufferIn(2193) when (flag_long='1') else '0';
	dataBufferOut(4552) <= dataBufferIn(2936) when (flag_long='1') else '0';
	dataBufferOut(4553) <= dataBufferIn(3679) when (flag_long='1') else '0';
	dataBufferOut(4554) <= dataBufferIn(4422) when (flag_long='1') else '0';
	dataBufferOut(4555) <= dataBufferIn(5165) when (flag_long='1') else '0';
	dataBufferOut(4556) <= dataBufferIn(5908) when (flag_long='1') else '0';
	dataBufferOut(4557) <= dataBufferIn( 507) when (flag_long='1') else '0';
	dataBufferOut(4558) <= dataBufferIn(1250) when (flag_long='1') else '0';
	dataBufferOut(4559) <= dataBufferIn(1993) when (flag_long='1') else '0';
	dataBufferOut(4560) <= dataBufferIn(2736) when (flag_long='1') else '0';
	dataBufferOut(4561) <= dataBufferIn(3479) when (flag_long='1') else '0';
	dataBufferOut(4562) <= dataBufferIn(4222) when (flag_long='1') else '0';
	dataBufferOut(4563) <= dataBufferIn(4965) when (flag_long='1') else '0';
	dataBufferOut(4564) <= dataBufferIn(5708) when (flag_long='1') else '0';
	dataBufferOut(4565) <= dataBufferIn( 307) when (flag_long='1') else '0';
	dataBufferOut(4566) <= dataBufferIn(1050) when (flag_long='1') else '0';
	dataBufferOut(4567) <= dataBufferIn(1793) when (flag_long='1') else '0';
	dataBufferOut(4568) <= dataBufferIn(2536) when (flag_long='1') else '0';
	dataBufferOut(4569) <= dataBufferIn(3279) when (flag_long='1') else '0';
	dataBufferOut(4570) <= dataBufferIn(4022) when (flag_long='1') else '0';
	dataBufferOut(4571) <= dataBufferIn(4765) when (flag_long='1') else '0';
	dataBufferOut(4572) <= dataBufferIn(5508) when (flag_long='1') else '0';
	dataBufferOut(4573) <= dataBufferIn( 107) when (flag_long='1') else '0';
	dataBufferOut(4574) <= dataBufferIn( 850) when (flag_long='1') else '0';
	dataBufferOut(4575) <= dataBufferIn(1593) when (flag_long='1') else '0';
	dataBufferOut(4576) <= dataBufferIn(2336) when (flag_long='1') else '0';
	dataBufferOut(4577) <= dataBufferIn(3079) when (flag_long='1') else '0';
	dataBufferOut(4578) <= dataBufferIn(3822) when (flag_long='1') else '0';
	dataBufferOut(4579) <= dataBufferIn(4565) when (flag_long='1') else '0';
	dataBufferOut(4580) <= dataBufferIn(5308) when (flag_long='1') else '0';
	dataBufferOut(4581) <= dataBufferIn(6051) when (flag_long='1') else '0';
	dataBufferOut(4582) <= dataBufferIn( 650) when (flag_long='1') else '0';
	dataBufferOut(4583) <= dataBufferIn(1393) when (flag_long='1') else '0';
	dataBufferOut(4584) <= dataBufferIn(2136) when (flag_long='1') else '0';
	dataBufferOut(4585) <= dataBufferIn(2879) when (flag_long='1') else '0';
	dataBufferOut(4586) <= dataBufferIn(3622) when (flag_long='1') else '0';
	dataBufferOut(4587) <= dataBufferIn(4365) when (flag_long='1') else '0';
	dataBufferOut(4588) <= dataBufferIn(5108) when (flag_long='1') else '0';
	dataBufferOut(4589) <= dataBufferIn(5851) when (flag_long='1') else '0';
	dataBufferOut(4590) <= dataBufferIn( 450) when (flag_long='1') else '0';
	dataBufferOut(4591) <= dataBufferIn(1193) when (flag_long='1') else '0';
	dataBufferOut(4592) <= dataBufferIn(1936) when (flag_long='1') else '0';
	dataBufferOut(4593) <= dataBufferIn(2679) when (flag_long='1') else '0';
	dataBufferOut(4594) <= dataBufferIn(3422) when (flag_long='1') else '0';
	dataBufferOut(4595) <= dataBufferIn(4165) when (flag_long='1') else '0';
	dataBufferOut(4596) <= dataBufferIn(4908) when (flag_long='1') else '0';
	dataBufferOut(4597) <= dataBufferIn(5651) when (flag_long='1') else '0';
	dataBufferOut(4598) <= dataBufferIn( 250) when (flag_long='1') else '0';
	dataBufferOut(4599) <= dataBufferIn( 993) when (flag_long='1') else '0';
	dataBufferOut(4600) <= dataBufferIn(1736) when (flag_long='1') else '0';
	dataBufferOut(4601) <= dataBufferIn(2479) when (flag_long='1') else '0';
	dataBufferOut(4602) <= dataBufferIn(3222) when (flag_long='1') else '0';
	dataBufferOut(4603) <= dataBufferIn(3965) when (flag_long='1') else '0';
	dataBufferOut(4604) <= dataBufferIn(4708) when (flag_long='1') else '0';
	dataBufferOut(4605) <= dataBufferIn(5451) when (flag_long='1') else '0';
	dataBufferOut(4606) <= dataBufferIn(  50) when (flag_long='1') else '0';
	dataBufferOut(4607) <= dataBufferIn( 793) when (flag_long='1') else '0';
	dataBufferOut(4608) <= dataBufferIn(1536) when (flag_long='1') else '0';
	dataBufferOut(4609) <= dataBufferIn(2279) when (flag_long='1') else '0';
	dataBufferOut(4610) <= dataBufferIn(3022) when (flag_long='1') else '0';
	dataBufferOut(4611) <= dataBufferIn(3765) when (flag_long='1') else '0';
	dataBufferOut(4612) <= dataBufferIn(4508) when (flag_long='1') else '0';
	dataBufferOut(4613) <= dataBufferIn(5251) when (flag_long='1') else '0';
	dataBufferOut(4614) <= dataBufferIn(5994) when (flag_long='1') else '0';
	dataBufferOut(4615) <= dataBufferIn( 593) when (flag_long='1') else '0';
	dataBufferOut(4616) <= dataBufferIn(1336) when (flag_long='1') else '0';
	dataBufferOut(4617) <= dataBufferIn(2079) when (flag_long='1') else '0';
	dataBufferOut(4618) <= dataBufferIn(2822) when (flag_long='1') else '0';
	dataBufferOut(4619) <= dataBufferIn(3565) when (flag_long='1') else '0';
	dataBufferOut(4620) <= dataBufferIn(4308) when (flag_long='1') else '0';
	dataBufferOut(4621) <= dataBufferIn(5051) when (flag_long='1') else '0';
	dataBufferOut(4622) <= dataBufferIn(5794) when (flag_long='1') else '0';
	dataBufferOut(4623) <= dataBufferIn( 393) when (flag_long='1') else '0';
	dataBufferOut(4624) <= dataBufferIn(1136) when (flag_long='1') else '0';
	dataBufferOut(4625) <= dataBufferIn(1879) when (flag_long='1') else '0';
	dataBufferOut(4626) <= dataBufferIn(2622) when (flag_long='1') else '0';
	dataBufferOut(4627) <= dataBufferIn(3365) when (flag_long='1') else '0';
	dataBufferOut(4628) <= dataBufferIn(4108) when (flag_long='1') else '0';
	dataBufferOut(4629) <= dataBufferIn(4851) when (flag_long='1') else '0';
	dataBufferOut(4630) <= dataBufferIn(5594) when (flag_long='1') else '0';
	dataBufferOut(4631) <= dataBufferIn( 193) when (flag_long='1') else '0';
	dataBufferOut(4632) <= dataBufferIn( 936) when (flag_long='1') else '0';
	dataBufferOut(4633) <= dataBufferIn(1679) when (flag_long='1') else '0';
	dataBufferOut(4634) <= dataBufferIn(2422) when (flag_long='1') else '0';
	dataBufferOut(4635) <= dataBufferIn(3165) when (flag_long='1') else '0';
	dataBufferOut(4636) <= dataBufferIn(3908) when (flag_long='1') else '0';
	dataBufferOut(4637) <= dataBufferIn(4651) when (flag_long='1') else '0';
	dataBufferOut(4638) <= dataBufferIn(5394) when (flag_long='1') else '0';
	dataBufferOut(4639) <= dataBufferIn(6137) when (flag_long='1') else '0';
	dataBufferOut(4640) <= dataBufferIn( 736) when (flag_long='1') else '0';
	dataBufferOut(4641) <= dataBufferIn(1479) when (flag_long='1') else '0';
	dataBufferOut(4642) <= dataBufferIn(2222) when (flag_long='1') else '0';
	dataBufferOut(4643) <= dataBufferIn(2965) when (flag_long='1') else '0';
	dataBufferOut(4644) <= dataBufferIn(3708) when (flag_long='1') else '0';
	dataBufferOut(4645) <= dataBufferIn(4451) when (flag_long='1') else '0';
	dataBufferOut(4646) <= dataBufferIn(5194) when (flag_long='1') else '0';
	dataBufferOut(4647) <= dataBufferIn(5937) when (flag_long='1') else '0';
	dataBufferOut(4648) <= dataBufferIn( 536) when (flag_long='1') else '0';
	dataBufferOut(4649) <= dataBufferIn(1279) when (flag_long='1') else '0';
	dataBufferOut(4650) <= dataBufferIn(2022) when (flag_long='1') else '0';
	dataBufferOut(4651) <= dataBufferIn(2765) when (flag_long='1') else '0';
	dataBufferOut(4652) <= dataBufferIn(3508) when (flag_long='1') else '0';
	dataBufferOut(4653) <= dataBufferIn(4251) when (flag_long='1') else '0';
	dataBufferOut(4654) <= dataBufferIn(4994) when (flag_long='1') else '0';
	dataBufferOut(4655) <= dataBufferIn(5737) when (flag_long='1') else '0';
	dataBufferOut(4656) <= dataBufferIn( 336) when (flag_long='1') else '0';
	dataBufferOut(4657) <= dataBufferIn(1079) when (flag_long='1') else '0';
	dataBufferOut(4658) <= dataBufferIn(1822) when (flag_long='1') else '0';
	dataBufferOut(4659) <= dataBufferIn(2565) when (flag_long='1') else '0';
	dataBufferOut(4660) <= dataBufferIn(3308) when (flag_long='1') else '0';
	dataBufferOut(4661) <= dataBufferIn(4051) when (flag_long='1') else '0';
	dataBufferOut(4662) <= dataBufferIn(4794) when (flag_long='1') else '0';
	dataBufferOut(4663) <= dataBufferIn(5537) when (flag_long='1') else '0';
	dataBufferOut(4664) <= dataBufferIn( 136) when (flag_long='1') else '0';
	dataBufferOut(4665) <= dataBufferIn( 879) when (flag_long='1') else '0';
	dataBufferOut(4666) <= dataBufferIn(1622) when (flag_long='1') else '0';
	dataBufferOut(4667) <= dataBufferIn(2365) when (flag_long='1') else '0';
	dataBufferOut(4668) <= dataBufferIn(3108) when (flag_long='1') else '0';
	dataBufferOut(4669) <= dataBufferIn(3851) when (flag_long='1') else '0';
	dataBufferOut(4670) <= dataBufferIn(4594) when (flag_long='1') else '0';
	dataBufferOut(4671) <= dataBufferIn(5337) when (flag_long='1') else '0';
	dataBufferOut(4672) <= dataBufferIn(6080) when (flag_long='1') else '0';
	dataBufferOut(4673) <= dataBufferIn( 679) when (flag_long='1') else '0';
	dataBufferOut(4674) <= dataBufferIn(1422) when (flag_long='1') else '0';
	dataBufferOut(4675) <= dataBufferIn(2165) when (flag_long='1') else '0';
	dataBufferOut(4676) <= dataBufferIn(2908) when (flag_long='1') else '0';
	dataBufferOut(4677) <= dataBufferIn(3651) when (flag_long='1') else '0';
	dataBufferOut(4678) <= dataBufferIn(4394) when (flag_long='1') else '0';
	dataBufferOut(4679) <= dataBufferIn(5137) when (flag_long='1') else '0';
	dataBufferOut(4680) <= dataBufferIn(5880) when (flag_long='1') else '0';
	dataBufferOut(4681) <= dataBufferIn( 479) when (flag_long='1') else '0';
	dataBufferOut(4682) <= dataBufferIn(1222) when (flag_long='1') else '0';
	dataBufferOut(4683) <= dataBufferIn(1965) when (flag_long='1') else '0';
	dataBufferOut(4684) <= dataBufferIn(2708) when (flag_long='1') else '0';
	dataBufferOut(4685) <= dataBufferIn(3451) when (flag_long='1') else '0';
	dataBufferOut(4686) <= dataBufferIn(4194) when (flag_long='1') else '0';
	dataBufferOut(4687) <= dataBufferIn(4937) when (flag_long='1') else '0';
	dataBufferOut(4688) <= dataBufferIn(5680) when (flag_long='1') else '0';
	dataBufferOut(4689) <= dataBufferIn( 279) when (flag_long='1') else '0';
	dataBufferOut(4690) <= dataBufferIn(1022) when (flag_long='1') else '0';
	dataBufferOut(4691) <= dataBufferIn(1765) when (flag_long='1') else '0';
	dataBufferOut(4692) <= dataBufferIn(2508) when (flag_long='1') else '0';
	dataBufferOut(4693) <= dataBufferIn(3251) when (flag_long='1') else '0';
	dataBufferOut(4694) <= dataBufferIn(3994) when (flag_long='1') else '0';
	dataBufferOut(4695) <= dataBufferIn(4737) when (flag_long='1') else '0';
	dataBufferOut(4696) <= dataBufferIn(5480) when (flag_long='1') else '0';
	dataBufferOut(4697) <= dataBufferIn(  79) when (flag_long='1') else '0';
	dataBufferOut(4698) <= dataBufferIn( 822) when (flag_long='1') else '0';
	dataBufferOut(4699) <= dataBufferIn(1565) when (flag_long='1') else '0';
	dataBufferOut(4700) <= dataBufferIn(2308) when (flag_long='1') else '0';
	dataBufferOut(4701) <= dataBufferIn(3051) when (flag_long='1') else '0';
	dataBufferOut(4702) <= dataBufferIn(3794) when (flag_long='1') else '0';
	dataBufferOut(4703) <= dataBufferIn(4537) when (flag_long='1') else '0';
	dataBufferOut(4704) <= dataBufferIn(5280) when (flag_long='1') else '0';
	dataBufferOut(4705) <= dataBufferIn(6023) when (flag_long='1') else '0';
	dataBufferOut(4706) <= dataBufferIn( 622) when (flag_long='1') else '0';
	dataBufferOut(4707) <= dataBufferIn(1365) when (flag_long='1') else '0';
	dataBufferOut(4708) <= dataBufferIn(2108) when (flag_long='1') else '0';
	dataBufferOut(4709) <= dataBufferIn(2851) when (flag_long='1') else '0';
	dataBufferOut(4710) <= dataBufferIn(3594) when (flag_long='1') else '0';
	dataBufferOut(4711) <= dataBufferIn(4337) when (flag_long='1') else '0';
	dataBufferOut(4712) <= dataBufferIn(5080) when (flag_long='1') else '0';
	dataBufferOut(4713) <= dataBufferIn(5823) when (flag_long='1') else '0';
	dataBufferOut(4714) <= dataBufferIn( 422) when (flag_long='1') else '0';
	dataBufferOut(4715) <= dataBufferIn(1165) when (flag_long='1') else '0';
	dataBufferOut(4716) <= dataBufferIn(1908) when (flag_long='1') else '0';
	dataBufferOut(4717) <= dataBufferIn(2651) when (flag_long='1') else '0';
	dataBufferOut(4718) <= dataBufferIn(3394) when (flag_long='1') else '0';
	dataBufferOut(4719) <= dataBufferIn(4137) when (flag_long='1') else '0';
	dataBufferOut(4720) <= dataBufferIn(4880) when (flag_long='1') else '0';
	dataBufferOut(4721) <= dataBufferIn(5623) when (flag_long='1') else '0';
	dataBufferOut(4722) <= dataBufferIn( 222) when (flag_long='1') else '0';
	dataBufferOut(4723) <= dataBufferIn( 965) when (flag_long='1') else '0';
	dataBufferOut(4724) <= dataBufferIn(1708) when (flag_long='1') else '0';
	dataBufferOut(4725) <= dataBufferIn(2451) when (flag_long='1') else '0';
	dataBufferOut(4726) <= dataBufferIn(3194) when (flag_long='1') else '0';
	dataBufferOut(4727) <= dataBufferIn(3937) when (flag_long='1') else '0';
	dataBufferOut(4728) <= dataBufferIn(4680) when (flag_long='1') else '0';
	dataBufferOut(4729) <= dataBufferIn(5423) when (flag_long='1') else '0';
	dataBufferOut(4730) <= dataBufferIn(  22) when (flag_long='1') else '0';
	dataBufferOut(4731) <= dataBufferIn( 765) when (flag_long='1') else '0';
	dataBufferOut(4732) <= dataBufferIn(1508) when (flag_long='1') else '0';
	dataBufferOut(4733) <= dataBufferIn(2251) when (flag_long='1') else '0';
	dataBufferOut(4734) <= dataBufferIn(2994) when (flag_long='1') else '0';
	dataBufferOut(4735) <= dataBufferIn(3737) when (flag_long='1') else '0';
	dataBufferOut(4736) <= dataBufferIn(4480) when (flag_long='1') else '0';
	dataBufferOut(4737) <= dataBufferIn(5223) when (flag_long='1') else '0';
	dataBufferOut(4738) <= dataBufferIn(5966) when (flag_long='1') else '0';
	dataBufferOut(4739) <= dataBufferIn( 565) when (flag_long='1') else '0';
	dataBufferOut(4740) <= dataBufferIn(1308) when (flag_long='1') else '0';
	dataBufferOut(4741) <= dataBufferIn(2051) when (flag_long='1') else '0';
	dataBufferOut(4742) <= dataBufferIn(2794) when (flag_long='1') else '0';
	dataBufferOut(4743) <= dataBufferIn(3537) when (flag_long='1') else '0';
	dataBufferOut(4744) <= dataBufferIn(4280) when (flag_long='1') else '0';
	dataBufferOut(4745) <= dataBufferIn(5023) when (flag_long='1') else '0';
	dataBufferOut(4746) <= dataBufferIn(5766) when (flag_long='1') else '0';
	dataBufferOut(4747) <= dataBufferIn( 365) when (flag_long='1') else '0';
	dataBufferOut(4748) <= dataBufferIn(1108) when (flag_long='1') else '0';
	dataBufferOut(4749) <= dataBufferIn(1851) when (flag_long='1') else '0';
	dataBufferOut(4750) <= dataBufferIn(2594) when (flag_long='1') else '0';
	dataBufferOut(4751) <= dataBufferIn(3337) when (flag_long='1') else '0';
	dataBufferOut(4752) <= dataBufferIn(4080) when (flag_long='1') else '0';
	dataBufferOut(4753) <= dataBufferIn(4823) when (flag_long='1') else '0';
	dataBufferOut(4754) <= dataBufferIn(5566) when (flag_long='1') else '0';
	dataBufferOut(4755) <= dataBufferIn( 165) when (flag_long='1') else '0';
	dataBufferOut(4756) <= dataBufferIn( 908) when (flag_long='1') else '0';
	dataBufferOut(4757) <= dataBufferIn(1651) when (flag_long='1') else '0';
	dataBufferOut(4758) <= dataBufferIn(2394) when (flag_long='1') else '0';
	dataBufferOut(4759) <= dataBufferIn(3137) when (flag_long='1') else '0';
	dataBufferOut(4760) <= dataBufferIn(3880) when (flag_long='1') else '0';
	dataBufferOut(4761) <= dataBufferIn(4623) when (flag_long='1') else '0';
	dataBufferOut(4762) <= dataBufferIn(5366) when (flag_long='1') else '0';
	dataBufferOut(4763) <= dataBufferIn(6109) when (flag_long='1') else '0';
	dataBufferOut(4764) <= dataBufferIn( 708) when (flag_long='1') else '0';
	dataBufferOut(4765) <= dataBufferIn(1451) when (flag_long='1') else '0';
	dataBufferOut(4766) <= dataBufferIn(2194) when (flag_long='1') else '0';
	dataBufferOut(4767) <= dataBufferIn(2937) when (flag_long='1') else '0';
	dataBufferOut(4768) <= dataBufferIn(3680) when (flag_long='1') else '0';
	dataBufferOut(4769) <= dataBufferIn(4423) when (flag_long='1') else '0';
	dataBufferOut(4770) <= dataBufferIn(5166) when (flag_long='1') else '0';
	dataBufferOut(4771) <= dataBufferIn(5909) when (flag_long='1') else '0';
	dataBufferOut(4772) <= dataBufferIn( 508) when (flag_long='1') else '0';
	dataBufferOut(4773) <= dataBufferIn(1251) when (flag_long='1') else '0';
	dataBufferOut(4774) <= dataBufferIn(1994) when (flag_long='1') else '0';
	dataBufferOut(4775) <= dataBufferIn(2737) when (flag_long='1') else '0';
	dataBufferOut(4776) <= dataBufferIn(3480) when (flag_long='1') else '0';
	dataBufferOut(4777) <= dataBufferIn(4223) when (flag_long='1') else '0';
	dataBufferOut(4778) <= dataBufferIn(4966) when (flag_long='1') else '0';
	dataBufferOut(4779) <= dataBufferIn(5709) when (flag_long='1') else '0';
	dataBufferOut(4780) <= dataBufferIn( 308) when (flag_long='1') else '0';
	dataBufferOut(4781) <= dataBufferIn(1051) when (flag_long='1') else '0';
	dataBufferOut(4782) <= dataBufferIn(1794) when (flag_long='1') else '0';
	dataBufferOut(4783) <= dataBufferIn(2537) when (flag_long='1') else '0';
	dataBufferOut(4784) <= dataBufferIn(3280) when (flag_long='1') else '0';
	dataBufferOut(4785) <= dataBufferIn(4023) when (flag_long='1') else '0';
	dataBufferOut(4786) <= dataBufferIn(4766) when (flag_long='1') else '0';
	dataBufferOut(4787) <= dataBufferIn(5509) when (flag_long='1') else '0';
	dataBufferOut(4788) <= dataBufferIn( 108) when (flag_long='1') else '0';
	dataBufferOut(4789) <= dataBufferIn( 851) when (flag_long='1') else '0';
	dataBufferOut(4790) <= dataBufferIn(1594) when (flag_long='1') else '0';
	dataBufferOut(4791) <= dataBufferIn(2337) when (flag_long='1') else '0';
	dataBufferOut(4792) <= dataBufferIn(3080) when (flag_long='1') else '0';
	dataBufferOut(4793) <= dataBufferIn(3823) when (flag_long='1') else '0';
	dataBufferOut(4794) <= dataBufferIn(4566) when (flag_long='1') else '0';
	dataBufferOut(4795) <= dataBufferIn(5309) when (flag_long='1') else '0';
	dataBufferOut(4796) <= dataBufferIn(6052) when (flag_long='1') else '0';
	dataBufferOut(4797) <= dataBufferIn( 651) when (flag_long='1') else '0';
	dataBufferOut(4798) <= dataBufferIn(1394) when (flag_long='1') else '0';
	dataBufferOut(4799) <= dataBufferIn(2137) when (flag_long='1') else '0';
	dataBufferOut(4800) <= dataBufferIn(2880) when (flag_long='1') else '0';
	dataBufferOut(4801) <= dataBufferIn(3623) when (flag_long='1') else '0';
	dataBufferOut(4802) <= dataBufferIn(4366) when (flag_long='1') else '0';
	dataBufferOut(4803) <= dataBufferIn(5109) when (flag_long='1') else '0';
	dataBufferOut(4804) <= dataBufferIn(5852) when (flag_long='1') else '0';
	dataBufferOut(4805) <= dataBufferIn( 451) when (flag_long='1') else '0';
	dataBufferOut(4806) <= dataBufferIn(1194) when (flag_long='1') else '0';
	dataBufferOut(4807) <= dataBufferIn(1937) when (flag_long='1') else '0';
	dataBufferOut(4808) <= dataBufferIn(2680) when (flag_long='1') else '0';
	dataBufferOut(4809) <= dataBufferIn(3423) when (flag_long='1') else '0';
	dataBufferOut(4810) <= dataBufferIn(4166) when (flag_long='1') else '0';
	dataBufferOut(4811) <= dataBufferIn(4909) when (flag_long='1') else '0';
	dataBufferOut(4812) <= dataBufferIn(5652) when (flag_long='1') else '0';
	dataBufferOut(4813) <= dataBufferIn( 251) when (flag_long='1') else '0';
	dataBufferOut(4814) <= dataBufferIn( 994) when (flag_long='1') else '0';
	dataBufferOut(4815) <= dataBufferIn(1737) when (flag_long='1') else '0';
	dataBufferOut(4816) <= dataBufferIn(2480) when (flag_long='1') else '0';
	dataBufferOut(4817) <= dataBufferIn(3223) when (flag_long='1') else '0';
	dataBufferOut(4818) <= dataBufferIn(3966) when (flag_long='1') else '0';
	dataBufferOut(4819) <= dataBufferIn(4709) when (flag_long='1') else '0';
	dataBufferOut(4820) <= dataBufferIn(5452) when (flag_long='1') else '0';
	dataBufferOut(4821) <= dataBufferIn(  51) when (flag_long='1') else '0';
	dataBufferOut(4822) <= dataBufferIn( 794) when (flag_long='1') else '0';
	dataBufferOut(4823) <= dataBufferIn(1537) when (flag_long='1') else '0';
	dataBufferOut(4824) <= dataBufferIn(2280) when (flag_long='1') else '0';
	dataBufferOut(4825) <= dataBufferIn(3023) when (flag_long='1') else '0';
	dataBufferOut(4826) <= dataBufferIn(3766) when (flag_long='1') else '0';
	dataBufferOut(4827) <= dataBufferIn(4509) when (flag_long='1') else '0';
	dataBufferOut(4828) <= dataBufferIn(5252) when (flag_long='1') else '0';
	dataBufferOut(4829) <= dataBufferIn(5995) when (flag_long='1') else '0';
	dataBufferOut(4830) <= dataBufferIn( 594) when (flag_long='1') else '0';
	dataBufferOut(4831) <= dataBufferIn(1337) when (flag_long='1') else '0';
	dataBufferOut(4832) <= dataBufferIn(2080) when (flag_long='1') else '0';
	dataBufferOut(4833) <= dataBufferIn(2823) when (flag_long='1') else '0';
	dataBufferOut(4834) <= dataBufferIn(3566) when (flag_long='1') else '0';
	dataBufferOut(4835) <= dataBufferIn(4309) when (flag_long='1') else '0';
	dataBufferOut(4836) <= dataBufferIn(5052) when (flag_long='1') else '0';
	dataBufferOut(4837) <= dataBufferIn(5795) when (flag_long='1') else '0';
	dataBufferOut(4838) <= dataBufferIn( 394) when (flag_long='1') else '0';
	dataBufferOut(4839) <= dataBufferIn(1137) when (flag_long='1') else '0';
	dataBufferOut(4840) <= dataBufferIn(1880) when (flag_long='1') else '0';
	dataBufferOut(4841) <= dataBufferIn(2623) when (flag_long='1') else '0';
	dataBufferOut(4842) <= dataBufferIn(3366) when (flag_long='1') else '0';
	dataBufferOut(4843) <= dataBufferIn(4109) when (flag_long='1') else '0';
	dataBufferOut(4844) <= dataBufferIn(4852) when (flag_long='1') else '0';
	dataBufferOut(4845) <= dataBufferIn(5595) when (flag_long='1') else '0';
	dataBufferOut(4846) <= dataBufferIn( 194) when (flag_long='1') else '0';
	dataBufferOut(4847) <= dataBufferIn( 937) when (flag_long='1') else '0';
	dataBufferOut(4848) <= dataBufferIn(1680) when (flag_long='1') else '0';
	dataBufferOut(4849) <= dataBufferIn(2423) when (flag_long='1') else '0';
	dataBufferOut(4850) <= dataBufferIn(3166) when (flag_long='1') else '0';
	dataBufferOut(4851) <= dataBufferIn(3909) when (flag_long='1') else '0';
	dataBufferOut(4852) <= dataBufferIn(4652) when (flag_long='1') else '0';
	dataBufferOut(4853) <= dataBufferIn(5395) when (flag_long='1') else '0';
	dataBufferOut(4854) <= dataBufferIn(6138) when (flag_long='1') else '0';
	dataBufferOut(4855) <= dataBufferIn( 737) when (flag_long='1') else '0';
	dataBufferOut(4856) <= dataBufferIn(1480) when (flag_long='1') else '0';
	dataBufferOut(4857) <= dataBufferIn(2223) when (flag_long='1') else '0';
	dataBufferOut(4858) <= dataBufferIn(2966) when (flag_long='1') else '0';
	dataBufferOut(4859) <= dataBufferIn(3709) when (flag_long='1') else '0';
	dataBufferOut(4860) <= dataBufferIn(4452) when (flag_long='1') else '0';
	dataBufferOut(4861) <= dataBufferIn(5195) when (flag_long='1') else '0';
	dataBufferOut(4862) <= dataBufferIn(5938) when (flag_long='1') else '0';
	dataBufferOut(4863) <= dataBufferIn( 537) when (flag_long='1') else '0';
	dataBufferOut(4864) <= dataBufferIn(1280) when (flag_long='1') else '0';
	dataBufferOut(4865) <= dataBufferIn(2023) when (flag_long='1') else '0';
	dataBufferOut(4866) <= dataBufferIn(2766) when (flag_long='1') else '0';
	dataBufferOut(4867) <= dataBufferIn(3509) when (flag_long='1') else '0';
	dataBufferOut(4868) <= dataBufferIn(4252) when (flag_long='1') else '0';
	dataBufferOut(4869) <= dataBufferIn(4995) when (flag_long='1') else '0';
	dataBufferOut(4870) <= dataBufferIn(5738) when (flag_long='1') else '0';
	dataBufferOut(4871) <= dataBufferIn( 337) when (flag_long='1') else '0';
	dataBufferOut(4872) <= dataBufferIn(1080) when (flag_long='1') else '0';
	dataBufferOut(4873) <= dataBufferIn(1823) when (flag_long='1') else '0';
	dataBufferOut(4874) <= dataBufferIn(2566) when (flag_long='1') else '0';
	dataBufferOut(4875) <= dataBufferIn(3309) when (flag_long='1') else '0';
	dataBufferOut(4876) <= dataBufferIn(4052) when (flag_long='1') else '0';
	dataBufferOut(4877) <= dataBufferIn(4795) when (flag_long='1') else '0';
	dataBufferOut(4878) <= dataBufferIn(5538) when (flag_long='1') else '0';
	dataBufferOut(4879) <= dataBufferIn( 137) when (flag_long='1') else '0';
	dataBufferOut(4880) <= dataBufferIn( 880) when (flag_long='1') else '0';
	dataBufferOut(4881) <= dataBufferIn(1623) when (flag_long='1') else '0';
	dataBufferOut(4882) <= dataBufferIn(2366) when (flag_long='1') else '0';
	dataBufferOut(4883) <= dataBufferIn(3109) when (flag_long='1') else '0';
	dataBufferOut(4884) <= dataBufferIn(3852) when (flag_long='1') else '0';
	dataBufferOut(4885) <= dataBufferIn(4595) when (flag_long='1') else '0';
	dataBufferOut(4886) <= dataBufferIn(5338) when (flag_long='1') else '0';
	dataBufferOut(4887) <= dataBufferIn(6081) when (flag_long='1') else '0';
	dataBufferOut(4888) <= dataBufferIn( 680) when (flag_long='1') else '0';
	dataBufferOut(4889) <= dataBufferIn(1423) when (flag_long='1') else '0';
	dataBufferOut(4890) <= dataBufferIn(2166) when (flag_long='1') else '0';
	dataBufferOut(4891) <= dataBufferIn(2909) when (flag_long='1') else '0';
	dataBufferOut(4892) <= dataBufferIn(3652) when (flag_long='1') else '0';
	dataBufferOut(4893) <= dataBufferIn(4395) when (flag_long='1') else '0';
	dataBufferOut(4894) <= dataBufferIn(5138) when (flag_long='1') else '0';
	dataBufferOut(4895) <= dataBufferIn(5881) when (flag_long='1') else '0';
	dataBufferOut(4896) <= dataBufferIn( 480) when (flag_long='1') else '0';
	dataBufferOut(4897) <= dataBufferIn(1223) when (flag_long='1') else '0';
	dataBufferOut(4898) <= dataBufferIn(1966) when (flag_long='1') else '0';
	dataBufferOut(4899) <= dataBufferIn(2709) when (flag_long='1') else '0';
	dataBufferOut(4900) <= dataBufferIn(3452) when (flag_long='1') else '0';
	dataBufferOut(4901) <= dataBufferIn(4195) when (flag_long='1') else '0';
	dataBufferOut(4902) <= dataBufferIn(4938) when (flag_long='1') else '0';
	dataBufferOut(4903) <= dataBufferIn(5681) when (flag_long='1') else '0';
	dataBufferOut(4904) <= dataBufferIn( 280) when (flag_long='1') else '0';
	dataBufferOut(4905) <= dataBufferIn(1023) when (flag_long='1') else '0';
	dataBufferOut(4906) <= dataBufferIn(1766) when (flag_long='1') else '0';
	dataBufferOut(4907) <= dataBufferIn(2509) when (flag_long='1') else '0';
	dataBufferOut(4908) <= dataBufferIn(3252) when (flag_long='1') else '0';
	dataBufferOut(4909) <= dataBufferIn(3995) when (flag_long='1') else '0';
	dataBufferOut(4910) <= dataBufferIn(4738) when (flag_long='1') else '0';
	dataBufferOut(4911) <= dataBufferIn(5481) when (flag_long='1') else '0';
	dataBufferOut(4912) <= dataBufferIn(  80) when (flag_long='1') else '0';
	dataBufferOut(4913) <= dataBufferIn( 823) when (flag_long='1') else '0';
	dataBufferOut(4914) <= dataBufferIn(1566) when (flag_long='1') else '0';
	dataBufferOut(4915) <= dataBufferIn(2309) when (flag_long='1') else '0';
	dataBufferOut(4916) <= dataBufferIn(3052) when (flag_long='1') else '0';
	dataBufferOut(4917) <= dataBufferIn(3795) when (flag_long='1') else '0';
	dataBufferOut(4918) <= dataBufferIn(4538) when (flag_long='1') else '0';
	dataBufferOut(4919) <= dataBufferIn(5281) when (flag_long='1') else '0';
	dataBufferOut(4920) <= dataBufferIn(6024) when (flag_long='1') else '0';
	dataBufferOut(4921) <= dataBufferIn( 623) when (flag_long='1') else '0';
	dataBufferOut(4922) <= dataBufferIn(1366) when (flag_long='1') else '0';
	dataBufferOut(4923) <= dataBufferIn(2109) when (flag_long='1') else '0';
	dataBufferOut(4924) <= dataBufferIn(2852) when (flag_long='1') else '0';
	dataBufferOut(4925) <= dataBufferIn(3595) when (flag_long='1') else '0';
	dataBufferOut(4926) <= dataBufferIn(4338) when (flag_long='1') else '0';
	dataBufferOut(4927) <= dataBufferIn(5081) when (flag_long='1') else '0';
	dataBufferOut(4928) <= dataBufferIn(5824) when (flag_long='1') else '0';
	dataBufferOut(4929) <= dataBufferIn( 423) when (flag_long='1') else '0';
	dataBufferOut(4930) <= dataBufferIn(1166) when (flag_long='1') else '0';
	dataBufferOut(4931) <= dataBufferIn(1909) when (flag_long='1') else '0';
	dataBufferOut(4932) <= dataBufferIn(2652) when (flag_long='1') else '0';
	dataBufferOut(4933) <= dataBufferIn(3395) when (flag_long='1') else '0';
	dataBufferOut(4934) <= dataBufferIn(4138) when (flag_long='1') else '0';
	dataBufferOut(4935) <= dataBufferIn(4881) when (flag_long='1') else '0';
	dataBufferOut(4936) <= dataBufferIn(5624) when (flag_long='1') else '0';
	dataBufferOut(4937) <= dataBufferIn( 223) when (flag_long='1') else '0';
	dataBufferOut(4938) <= dataBufferIn( 966) when (flag_long='1') else '0';
	dataBufferOut(4939) <= dataBufferIn(1709) when (flag_long='1') else '0';
	dataBufferOut(4940) <= dataBufferIn(2452) when (flag_long='1') else '0';
	dataBufferOut(4941) <= dataBufferIn(3195) when (flag_long='1') else '0';
	dataBufferOut(4942) <= dataBufferIn(3938) when (flag_long='1') else '0';
	dataBufferOut(4943) <= dataBufferIn(4681) when (flag_long='1') else '0';
	dataBufferOut(4944) <= dataBufferIn(5424) when (flag_long='1') else '0';
	dataBufferOut(4945) <= dataBufferIn(  23) when (flag_long='1') else '0';
	dataBufferOut(4946) <= dataBufferIn( 766) when (flag_long='1') else '0';
	dataBufferOut(4947) <= dataBufferIn(1509) when (flag_long='1') else '0';
	dataBufferOut(4948) <= dataBufferIn(2252) when (flag_long='1') else '0';
	dataBufferOut(4949) <= dataBufferIn(2995) when (flag_long='1') else '0';
	dataBufferOut(4950) <= dataBufferIn(3738) when (flag_long='1') else '0';
	dataBufferOut(4951) <= dataBufferIn(4481) when (flag_long='1') else '0';
	dataBufferOut(4952) <= dataBufferIn(5224) when (flag_long='1') else '0';
	dataBufferOut(4953) <= dataBufferIn(5967) when (flag_long='1') else '0';
	dataBufferOut(4954) <= dataBufferIn( 566) when (flag_long='1') else '0';
	dataBufferOut(4955) <= dataBufferIn(1309) when (flag_long='1') else '0';
	dataBufferOut(4956) <= dataBufferIn(2052) when (flag_long='1') else '0';
	dataBufferOut(4957) <= dataBufferIn(2795) when (flag_long='1') else '0';
	dataBufferOut(4958) <= dataBufferIn(3538) when (flag_long='1') else '0';
	dataBufferOut(4959) <= dataBufferIn(4281) when (flag_long='1') else '0';
	dataBufferOut(4960) <= dataBufferIn(5024) when (flag_long='1') else '0';
	dataBufferOut(4961) <= dataBufferIn(5767) when (flag_long='1') else '0';
	dataBufferOut(4962) <= dataBufferIn( 366) when (flag_long='1') else '0';
	dataBufferOut(4963) <= dataBufferIn(1109) when (flag_long='1') else '0';
	dataBufferOut(4964) <= dataBufferIn(1852) when (flag_long='1') else '0';
	dataBufferOut(4965) <= dataBufferIn(2595) when (flag_long='1') else '0';
	dataBufferOut(4966) <= dataBufferIn(3338) when (flag_long='1') else '0';
	dataBufferOut(4967) <= dataBufferIn(4081) when (flag_long='1') else '0';
	dataBufferOut(4968) <= dataBufferIn(4824) when (flag_long='1') else '0';
	dataBufferOut(4969) <= dataBufferIn(5567) when (flag_long='1') else '0';
	dataBufferOut(4970) <= dataBufferIn( 166) when (flag_long='1') else '0';
	dataBufferOut(4971) <= dataBufferIn( 909) when (flag_long='1') else '0';
	dataBufferOut(4972) <= dataBufferIn(1652) when (flag_long='1') else '0';
	dataBufferOut(4973) <= dataBufferIn(2395) when (flag_long='1') else '0';
	dataBufferOut(4974) <= dataBufferIn(3138) when (flag_long='1') else '0';
	dataBufferOut(4975) <= dataBufferIn(3881) when (flag_long='1') else '0';
	dataBufferOut(4976) <= dataBufferIn(4624) when (flag_long='1') else '0';
	dataBufferOut(4977) <= dataBufferIn(5367) when (flag_long='1') else '0';
	dataBufferOut(4978) <= dataBufferIn(6110) when (flag_long='1') else '0';
	dataBufferOut(4979) <= dataBufferIn( 709) when (flag_long='1') else '0';
	dataBufferOut(4980) <= dataBufferIn(1452) when (flag_long='1') else '0';
	dataBufferOut(4981) <= dataBufferIn(2195) when (flag_long='1') else '0';
	dataBufferOut(4982) <= dataBufferIn(2938) when (flag_long='1') else '0';
	dataBufferOut(4983) <= dataBufferIn(3681) when (flag_long='1') else '0';
	dataBufferOut(4984) <= dataBufferIn(4424) when (flag_long='1') else '0';
	dataBufferOut(4985) <= dataBufferIn(5167) when (flag_long='1') else '0';
	dataBufferOut(4986) <= dataBufferIn(5910) when (flag_long='1') else '0';
	dataBufferOut(4987) <= dataBufferIn( 509) when (flag_long='1') else '0';
	dataBufferOut(4988) <= dataBufferIn(1252) when (flag_long='1') else '0';
	dataBufferOut(4989) <= dataBufferIn(1995) when (flag_long='1') else '0';
	dataBufferOut(4990) <= dataBufferIn(2738) when (flag_long='1') else '0';
	dataBufferOut(4991) <= dataBufferIn(3481) when (flag_long='1') else '0';
	dataBufferOut(4992) <= dataBufferIn(4224) when (flag_long='1') else '0';
	dataBufferOut(4993) <= dataBufferIn(4967) when (flag_long='1') else '0';
	dataBufferOut(4994) <= dataBufferIn(5710) when (flag_long='1') else '0';
	dataBufferOut(4995) <= dataBufferIn( 309) when (flag_long='1') else '0';
	dataBufferOut(4996) <= dataBufferIn(1052) when (flag_long='1') else '0';
	dataBufferOut(4997) <= dataBufferIn(1795) when (flag_long='1') else '0';
	dataBufferOut(4998) <= dataBufferIn(2538) when (flag_long='1') else '0';
	dataBufferOut(4999) <= dataBufferIn(3281) when (flag_long='1') else '0';
	dataBufferOut(5000) <= dataBufferIn(4024) when (flag_long='1') else '0';
	dataBufferOut(5001) <= dataBufferIn(4767) when (flag_long='1') else '0';
	dataBufferOut(5002) <= dataBufferIn(5510) when (flag_long='1') else '0';
	dataBufferOut(5003) <= dataBufferIn( 109) when (flag_long='1') else '0';
	dataBufferOut(5004) <= dataBufferIn( 852) when (flag_long='1') else '0';
	dataBufferOut(5005) <= dataBufferIn(1595) when (flag_long='1') else '0';
	dataBufferOut(5006) <= dataBufferIn(2338) when (flag_long='1') else '0';
	dataBufferOut(5007) <= dataBufferIn(3081) when (flag_long='1') else '0';
	dataBufferOut(5008) <= dataBufferIn(3824) when (flag_long='1') else '0';
	dataBufferOut(5009) <= dataBufferIn(4567) when (flag_long='1') else '0';
	dataBufferOut(5010) <= dataBufferIn(5310) when (flag_long='1') else '0';
	dataBufferOut(5011) <= dataBufferIn(6053) when (flag_long='1') else '0';
	dataBufferOut(5012) <= dataBufferIn( 652) when (flag_long='1') else '0';
	dataBufferOut(5013) <= dataBufferIn(1395) when (flag_long='1') else '0';
	dataBufferOut(5014) <= dataBufferIn(2138) when (flag_long='1') else '0';
	dataBufferOut(5015) <= dataBufferIn(2881) when (flag_long='1') else '0';
	dataBufferOut(5016) <= dataBufferIn(3624) when (flag_long='1') else '0';
	dataBufferOut(5017) <= dataBufferIn(4367) when (flag_long='1') else '0';
	dataBufferOut(5018) <= dataBufferIn(5110) when (flag_long='1') else '0';
	dataBufferOut(5019) <= dataBufferIn(5853) when (flag_long='1') else '0';
	dataBufferOut(5020) <= dataBufferIn( 452) when (flag_long='1') else '0';
	dataBufferOut(5021) <= dataBufferIn(1195) when (flag_long='1') else '0';
	dataBufferOut(5022) <= dataBufferIn(1938) when (flag_long='1') else '0';
	dataBufferOut(5023) <= dataBufferIn(2681) when (flag_long='1') else '0';
	dataBufferOut(5024) <= dataBufferIn(3424) when (flag_long='1') else '0';
	dataBufferOut(5025) <= dataBufferIn(4167) when (flag_long='1') else '0';
	dataBufferOut(5026) <= dataBufferIn(4910) when (flag_long='1') else '0';
	dataBufferOut(5027) <= dataBufferIn(5653) when (flag_long='1') else '0';
	dataBufferOut(5028) <= dataBufferIn( 252) when (flag_long='1') else '0';
	dataBufferOut(5029) <= dataBufferIn( 995) when (flag_long='1') else '0';
	dataBufferOut(5030) <= dataBufferIn(1738) when (flag_long='1') else '0';
	dataBufferOut(5031) <= dataBufferIn(2481) when (flag_long='1') else '0';
	dataBufferOut(5032) <= dataBufferIn(3224) when (flag_long='1') else '0';
	dataBufferOut(5033) <= dataBufferIn(3967) when (flag_long='1') else '0';
	dataBufferOut(5034) <= dataBufferIn(4710) when (flag_long='1') else '0';
	dataBufferOut(5035) <= dataBufferIn(5453) when (flag_long='1') else '0';
	dataBufferOut(5036) <= dataBufferIn(  52) when (flag_long='1') else '0';
	dataBufferOut(5037) <= dataBufferIn( 795) when (flag_long='1') else '0';
	dataBufferOut(5038) <= dataBufferIn(1538) when (flag_long='1') else '0';
	dataBufferOut(5039) <= dataBufferIn(2281) when (flag_long='1') else '0';
	dataBufferOut(5040) <= dataBufferIn(3024) when (flag_long='1') else '0';
	dataBufferOut(5041) <= dataBufferIn(3767) when (flag_long='1') else '0';
	dataBufferOut(5042) <= dataBufferIn(4510) when (flag_long='1') else '0';
	dataBufferOut(5043) <= dataBufferIn(5253) when (flag_long='1') else '0';
	dataBufferOut(5044) <= dataBufferIn(5996) when (flag_long='1') else '0';
	dataBufferOut(5045) <= dataBufferIn( 595) when (flag_long='1') else '0';
	dataBufferOut(5046) <= dataBufferIn(1338) when (flag_long='1') else '0';
	dataBufferOut(5047) <= dataBufferIn(2081) when (flag_long='1') else '0';
	dataBufferOut(5048) <= dataBufferIn(2824) when (flag_long='1') else '0';
	dataBufferOut(5049) <= dataBufferIn(3567) when (flag_long='1') else '0';
	dataBufferOut(5050) <= dataBufferIn(4310) when (flag_long='1') else '0';
	dataBufferOut(5051) <= dataBufferIn(5053) when (flag_long='1') else '0';
	dataBufferOut(5052) <= dataBufferIn(5796) when (flag_long='1') else '0';
	dataBufferOut(5053) <= dataBufferIn( 395) when (flag_long='1') else '0';
	dataBufferOut(5054) <= dataBufferIn(1138) when (flag_long='1') else '0';
	dataBufferOut(5055) <= dataBufferIn(1881) when (flag_long='1') else '0';
	dataBufferOut(5056) <= dataBufferIn(2624) when (flag_long='1') else '0';
	dataBufferOut(5057) <= dataBufferIn(3367) when (flag_long='1') else '0';
	dataBufferOut(5058) <= dataBufferIn(4110) when (flag_long='1') else '0';
	dataBufferOut(5059) <= dataBufferIn(4853) when (flag_long='1') else '0';
	dataBufferOut(5060) <= dataBufferIn(5596) when (flag_long='1') else '0';
	dataBufferOut(5061) <= dataBufferIn( 195) when (flag_long='1') else '0';
	dataBufferOut(5062) <= dataBufferIn( 938) when (flag_long='1') else '0';
	dataBufferOut(5063) <= dataBufferIn(1681) when (flag_long='1') else '0';
	dataBufferOut(5064) <= dataBufferIn(2424) when (flag_long='1') else '0';
	dataBufferOut(5065) <= dataBufferIn(3167) when (flag_long='1') else '0';
	dataBufferOut(5066) <= dataBufferIn(3910) when (flag_long='1') else '0';
	dataBufferOut(5067) <= dataBufferIn(4653) when (flag_long='1') else '0';
	dataBufferOut(5068) <= dataBufferIn(5396) when (flag_long='1') else '0';
	dataBufferOut(5069) <= dataBufferIn(6139) when (flag_long='1') else '0';
	dataBufferOut(5070) <= dataBufferIn( 738) when (flag_long='1') else '0';
	dataBufferOut(5071) <= dataBufferIn(1481) when (flag_long='1') else '0';
	dataBufferOut(5072) <= dataBufferIn(2224) when (flag_long='1') else '0';
	dataBufferOut(5073) <= dataBufferIn(2967) when (flag_long='1') else '0';
	dataBufferOut(5074) <= dataBufferIn(3710) when (flag_long='1') else '0';
	dataBufferOut(5075) <= dataBufferIn(4453) when (flag_long='1') else '0';
	dataBufferOut(5076) <= dataBufferIn(5196) when (flag_long='1') else '0';
	dataBufferOut(5077) <= dataBufferIn(5939) when (flag_long='1') else '0';
	dataBufferOut(5078) <= dataBufferIn( 538) when (flag_long='1') else '0';
	dataBufferOut(5079) <= dataBufferIn(1281) when (flag_long='1') else '0';
	dataBufferOut(5080) <= dataBufferIn(2024) when (flag_long='1') else '0';
	dataBufferOut(5081) <= dataBufferIn(2767) when (flag_long='1') else '0';
	dataBufferOut(5082) <= dataBufferIn(3510) when (flag_long='1') else '0';
	dataBufferOut(5083) <= dataBufferIn(4253) when (flag_long='1') else '0';
	dataBufferOut(5084) <= dataBufferIn(4996) when (flag_long='1') else '0';
	dataBufferOut(5085) <= dataBufferIn(5739) when (flag_long='1') else '0';
	dataBufferOut(5086) <= dataBufferIn( 338) when (flag_long='1') else '0';
	dataBufferOut(5087) <= dataBufferIn(1081) when (flag_long='1') else '0';
	dataBufferOut(5088) <= dataBufferIn(1824) when (flag_long='1') else dataBufferIn(5088);
	dataBufferOut(5089) <= dataBufferIn(2567) when (flag_long='1') else dataBufferIn(5171);
	dataBufferOut(5090) <= dataBufferIn(3310) when (flag_long='1') else dataBufferIn(5254);
	dataBufferOut(5091) <= dataBufferIn(4053) when (flag_long='1') else dataBufferIn(5337);
	dataBufferOut(5092) <= dataBufferIn(4796) when (flag_long='1') else dataBufferIn(5420);
	dataBufferOut(5093) <= dataBufferIn(5539) when (flag_long='1') else dataBufferIn(5503);
	dataBufferOut(5094) <= dataBufferIn( 138) when (flag_long='1') else dataBufferIn(5586);
	dataBufferOut(5095) <= dataBufferIn( 881) when (flag_long='1') else dataBufferIn(5669);
	dataBufferOut(5096) <= dataBufferIn(1624) when (flag_long='1') else dataBufferIn(5752);
	dataBufferOut(5097) <= dataBufferIn(2367) when (flag_long='1') else dataBufferIn(5835);
	dataBufferOut(5098) <= dataBufferIn(3110) when (flag_long='1') else dataBufferIn(5918);
	dataBufferOut(5099) <= dataBufferIn(3853) when (flag_long='1') else dataBufferIn(6001);
	dataBufferOut(5100) <= dataBufferIn(4596) when (flag_long='1') else dataBufferIn(6084);
	dataBufferOut(5101) <= dataBufferIn(5339) when (flag_long='1') else dataBufferIn(5111);
	dataBufferOut(5102) <= dataBufferIn(6082) when (flag_long='1') else dataBufferIn(5194);
	dataBufferOut(5103) <= dataBufferIn( 681) when (flag_long='1') else dataBufferIn(5277);
	dataBufferOut(5104) <= dataBufferIn(1424) when (flag_long='1') else dataBufferIn(5360);
	dataBufferOut(5105) <= dataBufferIn(2167) when (flag_long='1') else dataBufferIn(5443);
	dataBufferOut(5106) <= dataBufferIn(2910) when (flag_long='1') else dataBufferIn(5526);
	dataBufferOut(5107) <= dataBufferIn(3653) when (flag_long='1') else dataBufferIn(5609);
	dataBufferOut(5108) <= dataBufferIn(4396) when (flag_long='1') else dataBufferIn(5692);
	dataBufferOut(5109) <= dataBufferIn(5139) when (flag_long='1') else dataBufferIn(5775);
	dataBufferOut(5110) <= dataBufferIn(5882) when (flag_long='1') else dataBufferIn(5858);
	dataBufferOut(5111) <= dataBufferIn( 481) when (flag_long='1') else dataBufferIn(5941);
	dataBufferOut(5112) <= dataBufferIn(1224) when (flag_long='1') else dataBufferIn(6024);
	dataBufferOut(5113) <= dataBufferIn(1967) when (flag_long='1') else dataBufferIn(6107);
	dataBufferOut(5114) <= dataBufferIn(2710) when (flag_long='1') else dataBufferIn(5134);
	dataBufferOut(5115) <= dataBufferIn(3453) when (flag_long='1') else dataBufferIn(5217);
	dataBufferOut(5116) <= dataBufferIn(4196) when (flag_long='1') else dataBufferIn(5300);
	dataBufferOut(5117) <= dataBufferIn(4939) when (flag_long='1') else dataBufferIn(5383);
	dataBufferOut(5118) <= dataBufferIn(5682) when (flag_long='1') else dataBufferIn(5466);
	dataBufferOut(5119) <= dataBufferIn( 281) when (flag_long='1') else dataBufferIn(5549);
	dataBufferOut(5120) <= dataBufferIn(1024) when (flag_long='1') else dataBufferIn(5632);
	dataBufferOut(5121) <= dataBufferIn(1767) when (flag_long='1') else dataBufferIn(5715);
	dataBufferOut(5122) <= dataBufferIn(2510) when (flag_long='1') else dataBufferIn(5798);
	dataBufferOut(5123) <= dataBufferIn(3253) when (flag_long='1') else dataBufferIn(5881);
	dataBufferOut(5124) <= dataBufferIn(3996) when (flag_long='1') else dataBufferIn(5964);
	dataBufferOut(5125) <= dataBufferIn(4739) when (flag_long='1') else dataBufferIn(6047);
	dataBufferOut(5126) <= dataBufferIn(5482) when (flag_long='1') else dataBufferIn(6130);
	dataBufferOut(5127) <= dataBufferIn(  81) when (flag_long='1') else dataBufferIn(5157);
	dataBufferOut(5128) <= dataBufferIn( 824) when (flag_long='1') else dataBufferIn(5240);
	dataBufferOut(5129) <= dataBufferIn(1567) when (flag_long='1') else dataBufferIn(5323);
	dataBufferOut(5130) <= dataBufferIn(2310) when (flag_long='1') else dataBufferIn(5406);
	dataBufferOut(5131) <= dataBufferIn(3053) when (flag_long='1') else dataBufferIn(5489);
	dataBufferOut(5132) <= dataBufferIn(3796) when (flag_long='1') else dataBufferIn(5572);
	dataBufferOut(5133) <= dataBufferIn(4539) when (flag_long='1') else dataBufferIn(5655);
	dataBufferOut(5134) <= dataBufferIn(5282) when (flag_long='1') else dataBufferIn(5738);
	dataBufferOut(5135) <= dataBufferIn(6025) when (flag_long='1') else dataBufferIn(5821);
	dataBufferOut(5136) <= dataBufferIn( 624) when (flag_long='1') else dataBufferIn(5904);
	dataBufferOut(5137) <= dataBufferIn(1367) when (flag_long='1') else dataBufferIn(5987);
	dataBufferOut(5138) <= dataBufferIn(2110) when (flag_long='1') else dataBufferIn(6070);
	dataBufferOut(5139) <= dataBufferIn(2853) when (flag_long='1') else dataBufferIn(5097);
	dataBufferOut(5140) <= dataBufferIn(3596) when (flag_long='1') else dataBufferIn(5180);
	dataBufferOut(5141) <= dataBufferIn(4339) when (flag_long='1') else dataBufferIn(5263);
	dataBufferOut(5142) <= dataBufferIn(5082) when (flag_long='1') else dataBufferIn(5346);
	dataBufferOut(5143) <= dataBufferIn(5825) when (flag_long='1') else dataBufferIn(5429);
	dataBufferOut(5144) <= dataBufferIn( 424) when (flag_long='1') else dataBufferIn(5512);
	dataBufferOut(5145) <= dataBufferIn(1167) when (flag_long='1') else dataBufferIn(5595);
	dataBufferOut(5146) <= dataBufferIn(1910) when (flag_long='1') else dataBufferIn(5678);
	dataBufferOut(5147) <= dataBufferIn(2653) when (flag_long='1') else dataBufferIn(5761);
	dataBufferOut(5148) <= dataBufferIn(3396) when (flag_long='1') else dataBufferIn(5844);
	dataBufferOut(5149) <= dataBufferIn(4139) when (flag_long='1') else dataBufferIn(5927);
	dataBufferOut(5150) <= dataBufferIn(4882) when (flag_long='1') else dataBufferIn(6010);
	dataBufferOut(5151) <= dataBufferIn(5625) when (flag_long='1') else dataBufferIn(6093);
	dataBufferOut(5152) <= dataBufferIn( 224) when (flag_long='1') else dataBufferIn(5120);
	dataBufferOut(5153) <= dataBufferIn( 967) when (flag_long='1') else dataBufferIn(5203);
	dataBufferOut(5154) <= dataBufferIn(1710) when (flag_long='1') else dataBufferIn(5286);
	dataBufferOut(5155) <= dataBufferIn(2453) when (flag_long='1') else dataBufferIn(5369);
	dataBufferOut(5156) <= dataBufferIn(3196) when (flag_long='1') else dataBufferIn(5452);
	dataBufferOut(5157) <= dataBufferIn(3939) when (flag_long='1') else dataBufferIn(5535);
	dataBufferOut(5158) <= dataBufferIn(4682) when (flag_long='1') else dataBufferIn(5618);
	dataBufferOut(5159) <= dataBufferIn(5425) when (flag_long='1') else dataBufferIn(5701);
	dataBufferOut(5160) <= dataBufferIn(  24) when (flag_long='1') else dataBufferIn(5784);
	dataBufferOut(5161) <= dataBufferIn( 767) when (flag_long='1') else dataBufferIn(5867);
	dataBufferOut(5162) <= dataBufferIn(1510) when (flag_long='1') else dataBufferIn(5950);
	dataBufferOut(5163) <= dataBufferIn(2253) when (flag_long='1') else dataBufferIn(6033);
	dataBufferOut(5164) <= dataBufferIn(2996) when (flag_long='1') else dataBufferIn(6116);
	dataBufferOut(5165) <= dataBufferIn(3739) when (flag_long='1') else dataBufferIn(5143);
	dataBufferOut(5166) <= dataBufferIn(4482) when (flag_long='1') else dataBufferIn(5226);
	dataBufferOut(5167) <= dataBufferIn(5225) when (flag_long='1') else dataBufferIn(5309);
	dataBufferOut(5168) <= dataBufferIn(5968) when (flag_long='1') else dataBufferIn(5392);
	dataBufferOut(5169) <= dataBufferIn( 567) when (flag_long='1') else dataBufferIn(5475);
	dataBufferOut(5170) <= dataBufferIn(1310) when (flag_long='1') else dataBufferIn(5558);
	dataBufferOut(5171) <= dataBufferIn(2053) when (flag_long='1') else dataBufferIn(5641);
	dataBufferOut(5172) <= dataBufferIn(2796) when (flag_long='1') else dataBufferIn(5724);
	dataBufferOut(5173) <= dataBufferIn(3539) when (flag_long='1') else dataBufferIn(5807);
	dataBufferOut(5174) <= dataBufferIn(4282) when (flag_long='1') else dataBufferIn(5890);
	dataBufferOut(5175) <= dataBufferIn(5025) when (flag_long='1') else dataBufferIn(5973);
	dataBufferOut(5176) <= dataBufferIn(5768) when (flag_long='1') else dataBufferIn(6056);
	dataBufferOut(5177) <= dataBufferIn( 367) when (flag_long='1') else dataBufferIn(6139);
	dataBufferOut(5178) <= dataBufferIn(1110) when (flag_long='1') else dataBufferIn(5166);
	dataBufferOut(5179) <= dataBufferIn(1853) when (flag_long='1') else dataBufferIn(5249);
	dataBufferOut(5180) <= dataBufferIn(2596) when (flag_long='1') else dataBufferIn(5332);
	dataBufferOut(5181) <= dataBufferIn(3339) when (flag_long='1') else dataBufferIn(5415);
	dataBufferOut(5182) <= dataBufferIn(4082) when (flag_long='1') else dataBufferIn(5498);
	dataBufferOut(5183) <= dataBufferIn(4825) when (flag_long='1') else dataBufferIn(5581);
	dataBufferOut(5184) <= dataBufferIn(5568) when (flag_long='1') else dataBufferIn(5664);
	dataBufferOut(5185) <= dataBufferIn( 167) when (flag_long='1') else dataBufferIn(5747);
	dataBufferOut(5186) <= dataBufferIn( 910) when (flag_long='1') else dataBufferIn(5830);
	dataBufferOut(5187) <= dataBufferIn(1653) when (flag_long='1') else dataBufferIn(5913);
	dataBufferOut(5188) <= dataBufferIn(2396) when (flag_long='1') else dataBufferIn(5996);
	dataBufferOut(5189) <= dataBufferIn(3139) when (flag_long='1') else dataBufferIn(6079);
	dataBufferOut(5190) <= dataBufferIn(3882) when (flag_long='1') else dataBufferIn(5106);
	dataBufferOut(5191) <= dataBufferIn(4625) when (flag_long='1') else dataBufferIn(5189);
	dataBufferOut(5192) <= dataBufferIn(5368) when (flag_long='1') else dataBufferIn(5272);
	dataBufferOut(5193) <= dataBufferIn(6111) when (flag_long='1') else dataBufferIn(5355);
	dataBufferOut(5194) <= dataBufferIn( 710) when (flag_long='1') else dataBufferIn(5438);
	dataBufferOut(5195) <= dataBufferIn(1453) when (flag_long='1') else dataBufferIn(5521);
	dataBufferOut(5196) <= dataBufferIn(2196) when (flag_long='1') else dataBufferIn(5604);
	dataBufferOut(5197) <= dataBufferIn(2939) when (flag_long='1') else dataBufferIn(5687);
	dataBufferOut(5198) <= dataBufferIn(3682) when (flag_long='1') else dataBufferIn(5770);
	dataBufferOut(5199) <= dataBufferIn(4425) when (flag_long='1') else dataBufferIn(5853);
	dataBufferOut(5200) <= dataBufferIn(5168) when (flag_long='1') else dataBufferIn(5936);
	dataBufferOut(5201) <= dataBufferIn(5911) when (flag_long='1') else dataBufferIn(6019);
	dataBufferOut(5202) <= dataBufferIn( 510) when (flag_long='1') else dataBufferIn(6102);
	dataBufferOut(5203) <= dataBufferIn(1253) when (flag_long='1') else dataBufferIn(5129);
	dataBufferOut(5204) <= dataBufferIn(1996) when (flag_long='1') else dataBufferIn(5212);
	dataBufferOut(5205) <= dataBufferIn(2739) when (flag_long='1') else dataBufferIn(5295);
	dataBufferOut(5206) <= dataBufferIn(3482) when (flag_long='1') else dataBufferIn(5378);
	dataBufferOut(5207) <= dataBufferIn(4225) when (flag_long='1') else dataBufferIn(5461);
	dataBufferOut(5208) <= dataBufferIn(4968) when (flag_long='1') else dataBufferIn(5544);
	dataBufferOut(5209) <= dataBufferIn(5711) when (flag_long='1') else dataBufferIn(5627);
	dataBufferOut(5210) <= dataBufferIn( 310) when (flag_long='1') else dataBufferIn(5710);
	dataBufferOut(5211) <= dataBufferIn(1053) when (flag_long='1') else dataBufferIn(5793);
	dataBufferOut(5212) <= dataBufferIn(1796) when (flag_long='1') else dataBufferIn(5876);
	dataBufferOut(5213) <= dataBufferIn(2539) when (flag_long='1') else dataBufferIn(5959);
	dataBufferOut(5214) <= dataBufferIn(3282) when (flag_long='1') else dataBufferIn(6042);
	dataBufferOut(5215) <= dataBufferIn(4025) when (flag_long='1') else dataBufferIn(6125);
	dataBufferOut(5216) <= dataBufferIn(4768) when (flag_long='1') else dataBufferIn(5152);
	dataBufferOut(5217) <= dataBufferIn(5511) when (flag_long='1') else dataBufferIn(5235);
	dataBufferOut(5218) <= dataBufferIn( 110) when (flag_long='1') else dataBufferIn(5318);
	dataBufferOut(5219) <= dataBufferIn( 853) when (flag_long='1') else dataBufferIn(5401);
	dataBufferOut(5220) <= dataBufferIn(1596) when (flag_long='1') else dataBufferIn(5484);
	dataBufferOut(5221) <= dataBufferIn(2339) when (flag_long='1') else dataBufferIn(5567);
	dataBufferOut(5222) <= dataBufferIn(3082) when (flag_long='1') else dataBufferIn(5650);
	dataBufferOut(5223) <= dataBufferIn(3825) when (flag_long='1') else dataBufferIn(5733);
	dataBufferOut(5224) <= dataBufferIn(4568) when (flag_long='1') else dataBufferIn(5816);
	dataBufferOut(5225) <= dataBufferIn(5311) when (flag_long='1') else dataBufferIn(5899);
	dataBufferOut(5226) <= dataBufferIn(6054) when (flag_long='1') else dataBufferIn(5982);
	dataBufferOut(5227) <= dataBufferIn( 653) when (flag_long='1') else dataBufferIn(6065);
	dataBufferOut(5228) <= dataBufferIn(1396) when (flag_long='1') else dataBufferIn(5092);
	dataBufferOut(5229) <= dataBufferIn(2139) when (flag_long='1') else dataBufferIn(5175);
	dataBufferOut(5230) <= dataBufferIn(2882) when (flag_long='1') else dataBufferIn(5258);
	dataBufferOut(5231) <= dataBufferIn(3625) when (flag_long='1') else dataBufferIn(5341);
	dataBufferOut(5232) <= dataBufferIn(4368) when (flag_long='1') else dataBufferIn(5424);
	dataBufferOut(5233) <= dataBufferIn(5111) when (flag_long='1') else dataBufferIn(5507);
	dataBufferOut(5234) <= dataBufferIn(5854) when (flag_long='1') else dataBufferIn(5590);
	dataBufferOut(5235) <= dataBufferIn( 453) when (flag_long='1') else dataBufferIn(5673);
	dataBufferOut(5236) <= dataBufferIn(1196) when (flag_long='1') else dataBufferIn(5756);
	dataBufferOut(5237) <= dataBufferIn(1939) when (flag_long='1') else dataBufferIn(5839);
	dataBufferOut(5238) <= dataBufferIn(2682) when (flag_long='1') else dataBufferIn(5922);
	dataBufferOut(5239) <= dataBufferIn(3425) when (flag_long='1') else dataBufferIn(6005);
	dataBufferOut(5240) <= dataBufferIn(4168) when (flag_long='1') else dataBufferIn(6088);
	dataBufferOut(5241) <= dataBufferIn(4911) when (flag_long='1') else dataBufferIn(5115);
	dataBufferOut(5242) <= dataBufferIn(5654) when (flag_long='1') else dataBufferIn(5198);
	dataBufferOut(5243) <= dataBufferIn( 253) when (flag_long='1') else dataBufferIn(5281);
	dataBufferOut(5244) <= dataBufferIn( 996) when (flag_long='1') else dataBufferIn(5364);
	dataBufferOut(5245) <= dataBufferIn(1739) when (flag_long='1') else dataBufferIn(5447);
	dataBufferOut(5246) <= dataBufferIn(2482) when (flag_long='1') else dataBufferIn(5530);
	dataBufferOut(5247) <= dataBufferIn(3225) when (flag_long='1') else dataBufferIn(5613);
	dataBufferOut(5248) <= dataBufferIn(3968) when (flag_long='1') else dataBufferIn(5696);
	dataBufferOut(5249) <= dataBufferIn(4711) when (flag_long='1') else dataBufferIn(5779);
	dataBufferOut(5250) <= dataBufferIn(5454) when (flag_long='1') else dataBufferIn(5862);
	dataBufferOut(5251) <= dataBufferIn(  53) when (flag_long='1') else dataBufferIn(5945);
	dataBufferOut(5252) <= dataBufferIn( 796) when (flag_long='1') else dataBufferIn(6028);
	dataBufferOut(5253) <= dataBufferIn(1539) when (flag_long='1') else dataBufferIn(6111);
	dataBufferOut(5254) <= dataBufferIn(2282) when (flag_long='1') else dataBufferIn(5138);
	dataBufferOut(5255) <= dataBufferIn(3025) when (flag_long='1') else dataBufferIn(5221);
	dataBufferOut(5256) <= dataBufferIn(3768) when (flag_long='1') else dataBufferIn(5304);
	dataBufferOut(5257) <= dataBufferIn(4511) when (flag_long='1') else dataBufferIn(5387);
	dataBufferOut(5258) <= dataBufferIn(5254) when (flag_long='1') else dataBufferIn(5470);
	dataBufferOut(5259) <= dataBufferIn(5997) when (flag_long='1') else dataBufferIn(5553);
	dataBufferOut(5260) <= dataBufferIn( 596) when (flag_long='1') else dataBufferIn(5636);
	dataBufferOut(5261) <= dataBufferIn(1339) when (flag_long='1') else dataBufferIn(5719);
	dataBufferOut(5262) <= dataBufferIn(2082) when (flag_long='1') else dataBufferIn(5802);
	dataBufferOut(5263) <= dataBufferIn(2825) when (flag_long='1') else dataBufferIn(5885);
	dataBufferOut(5264) <= dataBufferIn(3568) when (flag_long='1') else dataBufferIn(5968);
	dataBufferOut(5265) <= dataBufferIn(4311) when (flag_long='1') else dataBufferIn(6051);
	dataBufferOut(5266) <= dataBufferIn(5054) when (flag_long='1') else dataBufferIn(6134);
	dataBufferOut(5267) <= dataBufferIn(5797) when (flag_long='1') else dataBufferIn(5161);
	dataBufferOut(5268) <= dataBufferIn( 396) when (flag_long='1') else dataBufferIn(5244);
	dataBufferOut(5269) <= dataBufferIn(1139) when (flag_long='1') else dataBufferIn(5327);
	dataBufferOut(5270) <= dataBufferIn(1882) when (flag_long='1') else dataBufferIn(5410);
	dataBufferOut(5271) <= dataBufferIn(2625) when (flag_long='1') else dataBufferIn(5493);
	dataBufferOut(5272) <= dataBufferIn(3368) when (flag_long='1') else dataBufferIn(5576);
	dataBufferOut(5273) <= dataBufferIn(4111) when (flag_long='1') else dataBufferIn(5659);
	dataBufferOut(5274) <= dataBufferIn(4854) when (flag_long='1') else dataBufferIn(5742);
	dataBufferOut(5275) <= dataBufferIn(5597) when (flag_long='1') else dataBufferIn(5825);
	dataBufferOut(5276) <= dataBufferIn( 196) when (flag_long='1') else dataBufferIn(5908);
	dataBufferOut(5277) <= dataBufferIn( 939) when (flag_long='1') else dataBufferIn(5991);
	dataBufferOut(5278) <= dataBufferIn(1682) when (flag_long='1') else dataBufferIn(6074);
	dataBufferOut(5279) <= dataBufferIn(2425) when (flag_long='1') else dataBufferIn(5101);
	dataBufferOut(5280) <= dataBufferIn(3168) when (flag_long='1') else dataBufferIn(5184);
	dataBufferOut(5281) <= dataBufferIn(3911) when (flag_long='1') else dataBufferIn(5267);
	dataBufferOut(5282) <= dataBufferIn(4654) when (flag_long='1') else dataBufferIn(5350);
	dataBufferOut(5283) <= dataBufferIn(5397) when (flag_long='1') else dataBufferIn(5433);
	dataBufferOut(5284) <= dataBufferIn(6140) when (flag_long='1') else dataBufferIn(5516);
	dataBufferOut(5285) <= dataBufferIn( 739) when (flag_long='1') else dataBufferIn(5599);
	dataBufferOut(5286) <= dataBufferIn(1482) when (flag_long='1') else dataBufferIn(5682);
	dataBufferOut(5287) <= dataBufferIn(2225) when (flag_long='1') else dataBufferIn(5765);
	dataBufferOut(5288) <= dataBufferIn(2968) when (flag_long='1') else dataBufferIn(5848);
	dataBufferOut(5289) <= dataBufferIn(3711) when (flag_long='1') else dataBufferIn(5931);
	dataBufferOut(5290) <= dataBufferIn(4454) when (flag_long='1') else dataBufferIn(6014);
	dataBufferOut(5291) <= dataBufferIn(5197) when (flag_long='1') else dataBufferIn(6097);
	dataBufferOut(5292) <= dataBufferIn(5940) when (flag_long='1') else dataBufferIn(5124);
	dataBufferOut(5293) <= dataBufferIn( 539) when (flag_long='1') else dataBufferIn(5207);
	dataBufferOut(5294) <= dataBufferIn(1282) when (flag_long='1') else dataBufferIn(5290);
	dataBufferOut(5295) <= dataBufferIn(2025) when (flag_long='1') else dataBufferIn(5373);
	dataBufferOut(5296) <= dataBufferIn(2768) when (flag_long='1') else dataBufferIn(5456);
	dataBufferOut(5297) <= dataBufferIn(3511) when (flag_long='1') else dataBufferIn(5539);
	dataBufferOut(5298) <= dataBufferIn(4254) when (flag_long='1') else dataBufferIn(5622);
	dataBufferOut(5299) <= dataBufferIn(4997) when (flag_long='1') else dataBufferIn(5705);
	dataBufferOut(5300) <= dataBufferIn(5740) when (flag_long='1') else dataBufferIn(5788);
	dataBufferOut(5301) <= dataBufferIn( 339) when (flag_long='1') else dataBufferIn(5871);
	dataBufferOut(5302) <= dataBufferIn(1082) when (flag_long='1') else dataBufferIn(5954);
	dataBufferOut(5303) <= dataBufferIn(1825) when (flag_long='1') else dataBufferIn(6037);
	dataBufferOut(5304) <= dataBufferIn(2568) when (flag_long='1') else dataBufferIn(6120);
	dataBufferOut(5305) <= dataBufferIn(3311) when (flag_long='1') else dataBufferIn(5147);
	dataBufferOut(5306) <= dataBufferIn(4054) when (flag_long='1') else dataBufferIn(5230);
	dataBufferOut(5307) <= dataBufferIn(4797) when (flag_long='1') else dataBufferIn(5313);
	dataBufferOut(5308) <= dataBufferIn(5540) when (flag_long='1') else dataBufferIn(5396);
	dataBufferOut(5309) <= dataBufferIn( 139) when (flag_long='1') else dataBufferIn(5479);
	dataBufferOut(5310) <= dataBufferIn( 882) when (flag_long='1') else dataBufferIn(5562);
	dataBufferOut(5311) <= dataBufferIn(1625) when (flag_long='1') else dataBufferIn(5645);
	dataBufferOut(5312) <= dataBufferIn(2368) when (flag_long='1') else dataBufferIn(5728);
	dataBufferOut(5313) <= dataBufferIn(3111) when (flag_long='1') else dataBufferIn(5811);
	dataBufferOut(5314) <= dataBufferIn(3854) when (flag_long='1') else dataBufferIn(5894);
	dataBufferOut(5315) <= dataBufferIn(4597) when (flag_long='1') else dataBufferIn(5977);
	dataBufferOut(5316) <= dataBufferIn(5340) when (flag_long='1') else dataBufferIn(6060);
	dataBufferOut(5317) <= dataBufferIn(6083) when (flag_long='1') else dataBufferIn(6143);
	dataBufferOut(5318) <= dataBufferIn( 682) when (flag_long='1') else dataBufferIn(5170);
	dataBufferOut(5319) <= dataBufferIn(1425) when (flag_long='1') else dataBufferIn(5253);
	dataBufferOut(5320) <= dataBufferIn(2168) when (flag_long='1') else dataBufferIn(5336);
	dataBufferOut(5321) <= dataBufferIn(2911) when (flag_long='1') else dataBufferIn(5419);
	dataBufferOut(5322) <= dataBufferIn(3654) when (flag_long='1') else dataBufferIn(5502);
	dataBufferOut(5323) <= dataBufferIn(4397) when (flag_long='1') else dataBufferIn(5585);
	dataBufferOut(5324) <= dataBufferIn(5140) when (flag_long='1') else dataBufferIn(5668);
	dataBufferOut(5325) <= dataBufferIn(5883) when (flag_long='1') else dataBufferIn(5751);
	dataBufferOut(5326) <= dataBufferIn( 482) when (flag_long='1') else dataBufferIn(5834);
	dataBufferOut(5327) <= dataBufferIn(1225) when (flag_long='1') else dataBufferIn(5917);
	dataBufferOut(5328) <= dataBufferIn(1968) when (flag_long='1') else dataBufferIn(6000);
	dataBufferOut(5329) <= dataBufferIn(2711) when (flag_long='1') else dataBufferIn(6083);
	dataBufferOut(5330) <= dataBufferIn(3454) when (flag_long='1') else dataBufferIn(5110);
	dataBufferOut(5331) <= dataBufferIn(4197) when (flag_long='1') else dataBufferIn(5193);
	dataBufferOut(5332) <= dataBufferIn(4940) when (flag_long='1') else dataBufferIn(5276);
	dataBufferOut(5333) <= dataBufferIn(5683) when (flag_long='1') else dataBufferIn(5359);
	dataBufferOut(5334) <= dataBufferIn( 282) when (flag_long='1') else dataBufferIn(5442);
	dataBufferOut(5335) <= dataBufferIn(1025) when (flag_long='1') else dataBufferIn(5525);
	dataBufferOut(5336) <= dataBufferIn(1768) when (flag_long='1') else dataBufferIn(5608);
	dataBufferOut(5337) <= dataBufferIn(2511) when (flag_long='1') else dataBufferIn(5691);
	dataBufferOut(5338) <= dataBufferIn(3254) when (flag_long='1') else dataBufferIn(5774);
	dataBufferOut(5339) <= dataBufferIn(3997) when (flag_long='1') else dataBufferIn(5857);
	dataBufferOut(5340) <= dataBufferIn(4740) when (flag_long='1') else dataBufferIn(5940);
	dataBufferOut(5341) <= dataBufferIn(5483) when (flag_long='1') else dataBufferIn(6023);
	dataBufferOut(5342) <= dataBufferIn(  82) when (flag_long='1') else dataBufferIn(6106);
	dataBufferOut(5343) <= dataBufferIn( 825) when (flag_long='1') else dataBufferIn(5133);
	dataBufferOut(5344) <= dataBufferIn(1568) when (flag_long='1') else dataBufferIn(5216);
	dataBufferOut(5345) <= dataBufferIn(2311) when (flag_long='1') else dataBufferIn(5299);
	dataBufferOut(5346) <= dataBufferIn(3054) when (flag_long='1') else dataBufferIn(5382);
	dataBufferOut(5347) <= dataBufferIn(3797) when (flag_long='1') else dataBufferIn(5465);
	dataBufferOut(5348) <= dataBufferIn(4540) when (flag_long='1') else dataBufferIn(5548);
	dataBufferOut(5349) <= dataBufferIn(5283) when (flag_long='1') else dataBufferIn(5631);
	dataBufferOut(5350) <= dataBufferIn(6026) when (flag_long='1') else dataBufferIn(5714);
	dataBufferOut(5351) <= dataBufferIn( 625) when (flag_long='1') else dataBufferIn(5797);
	dataBufferOut(5352) <= dataBufferIn(1368) when (flag_long='1') else dataBufferIn(5880);
	dataBufferOut(5353) <= dataBufferIn(2111) when (flag_long='1') else dataBufferIn(5963);
	dataBufferOut(5354) <= dataBufferIn(2854) when (flag_long='1') else dataBufferIn(6046);
	dataBufferOut(5355) <= dataBufferIn(3597) when (flag_long='1') else dataBufferIn(6129);
	dataBufferOut(5356) <= dataBufferIn(4340) when (flag_long='1') else dataBufferIn(5156);
	dataBufferOut(5357) <= dataBufferIn(5083) when (flag_long='1') else dataBufferIn(5239);
	dataBufferOut(5358) <= dataBufferIn(5826) when (flag_long='1') else dataBufferIn(5322);
	dataBufferOut(5359) <= dataBufferIn( 425) when (flag_long='1') else dataBufferIn(5405);
	dataBufferOut(5360) <= dataBufferIn(1168) when (flag_long='1') else dataBufferIn(5488);
	dataBufferOut(5361) <= dataBufferIn(1911) when (flag_long='1') else dataBufferIn(5571);
	dataBufferOut(5362) <= dataBufferIn(2654) when (flag_long='1') else dataBufferIn(5654);
	dataBufferOut(5363) <= dataBufferIn(3397) when (flag_long='1') else dataBufferIn(5737);
	dataBufferOut(5364) <= dataBufferIn(4140) when (flag_long='1') else dataBufferIn(5820);
	dataBufferOut(5365) <= dataBufferIn(4883) when (flag_long='1') else dataBufferIn(5903);
	dataBufferOut(5366) <= dataBufferIn(5626) when (flag_long='1') else dataBufferIn(5986);
	dataBufferOut(5367) <= dataBufferIn( 225) when (flag_long='1') else dataBufferIn(6069);
	dataBufferOut(5368) <= dataBufferIn( 968) when (flag_long='1') else dataBufferIn(5096);
	dataBufferOut(5369) <= dataBufferIn(1711) when (flag_long='1') else dataBufferIn(5179);
	dataBufferOut(5370) <= dataBufferIn(2454) when (flag_long='1') else dataBufferIn(5262);
	dataBufferOut(5371) <= dataBufferIn(3197) when (flag_long='1') else dataBufferIn(5345);
	dataBufferOut(5372) <= dataBufferIn(3940) when (flag_long='1') else dataBufferIn(5428);
	dataBufferOut(5373) <= dataBufferIn(4683) when (flag_long='1') else dataBufferIn(5511);
	dataBufferOut(5374) <= dataBufferIn(5426) when (flag_long='1') else dataBufferIn(5594);
	dataBufferOut(5375) <= dataBufferIn(  25) when (flag_long='1') else dataBufferIn(5677);
	dataBufferOut(5376) <= dataBufferIn( 768) when (flag_long='1') else dataBufferIn(5760);
	dataBufferOut(5377) <= dataBufferIn(1511) when (flag_long='1') else dataBufferIn(5843);
	dataBufferOut(5378) <= dataBufferIn(2254) when (flag_long='1') else dataBufferIn(5926);
	dataBufferOut(5379) <= dataBufferIn(2997) when (flag_long='1') else dataBufferIn(6009);
	dataBufferOut(5380) <= dataBufferIn(3740) when (flag_long='1') else dataBufferIn(6092);
	dataBufferOut(5381) <= dataBufferIn(4483) when (flag_long='1') else dataBufferIn(5119);
	dataBufferOut(5382) <= dataBufferIn(5226) when (flag_long='1') else dataBufferIn(5202);
	dataBufferOut(5383) <= dataBufferIn(5969) when (flag_long='1') else dataBufferIn(5285);
	dataBufferOut(5384) <= dataBufferIn( 568) when (flag_long='1') else dataBufferIn(5368);
	dataBufferOut(5385) <= dataBufferIn(1311) when (flag_long='1') else dataBufferIn(5451);
	dataBufferOut(5386) <= dataBufferIn(2054) when (flag_long='1') else dataBufferIn(5534);
	dataBufferOut(5387) <= dataBufferIn(2797) when (flag_long='1') else dataBufferIn(5617);
	dataBufferOut(5388) <= dataBufferIn(3540) when (flag_long='1') else dataBufferIn(5700);
	dataBufferOut(5389) <= dataBufferIn(4283) when (flag_long='1') else dataBufferIn(5783);
	dataBufferOut(5390) <= dataBufferIn(5026) when (flag_long='1') else dataBufferIn(5866);
	dataBufferOut(5391) <= dataBufferIn(5769) when (flag_long='1') else dataBufferIn(5949);
	dataBufferOut(5392) <= dataBufferIn( 368) when (flag_long='1') else dataBufferIn(6032);
	dataBufferOut(5393) <= dataBufferIn(1111) when (flag_long='1') else dataBufferIn(6115);
	dataBufferOut(5394) <= dataBufferIn(1854) when (flag_long='1') else dataBufferIn(5142);
	dataBufferOut(5395) <= dataBufferIn(2597) when (flag_long='1') else dataBufferIn(5225);
	dataBufferOut(5396) <= dataBufferIn(3340) when (flag_long='1') else dataBufferIn(5308);
	dataBufferOut(5397) <= dataBufferIn(4083) when (flag_long='1') else dataBufferIn(5391);
	dataBufferOut(5398) <= dataBufferIn(4826) when (flag_long='1') else dataBufferIn(5474);
	dataBufferOut(5399) <= dataBufferIn(5569) when (flag_long='1') else dataBufferIn(5557);
	dataBufferOut(5400) <= dataBufferIn( 168) when (flag_long='1') else dataBufferIn(5640);
	dataBufferOut(5401) <= dataBufferIn( 911) when (flag_long='1') else dataBufferIn(5723);
	dataBufferOut(5402) <= dataBufferIn(1654) when (flag_long='1') else dataBufferIn(5806);
	dataBufferOut(5403) <= dataBufferIn(2397) when (flag_long='1') else dataBufferIn(5889);
	dataBufferOut(5404) <= dataBufferIn(3140) when (flag_long='1') else dataBufferIn(5972);
	dataBufferOut(5405) <= dataBufferIn(3883) when (flag_long='1') else dataBufferIn(6055);
	dataBufferOut(5406) <= dataBufferIn(4626) when (flag_long='1') else dataBufferIn(6138);
	dataBufferOut(5407) <= dataBufferIn(5369) when (flag_long='1') else dataBufferIn(5165);
	dataBufferOut(5408) <= dataBufferIn(6112) when (flag_long='1') else dataBufferIn(5248);
	dataBufferOut(5409) <= dataBufferIn( 711) when (flag_long='1') else dataBufferIn(5331);
	dataBufferOut(5410) <= dataBufferIn(1454) when (flag_long='1') else dataBufferIn(5414);
	dataBufferOut(5411) <= dataBufferIn(2197) when (flag_long='1') else dataBufferIn(5497);
	dataBufferOut(5412) <= dataBufferIn(2940) when (flag_long='1') else dataBufferIn(5580);
	dataBufferOut(5413) <= dataBufferIn(3683) when (flag_long='1') else dataBufferIn(5663);
	dataBufferOut(5414) <= dataBufferIn(4426) when (flag_long='1') else dataBufferIn(5746);
	dataBufferOut(5415) <= dataBufferIn(5169) when (flag_long='1') else dataBufferIn(5829);
	dataBufferOut(5416) <= dataBufferIn(5912) when (flag_long='1') else dataBufferIn(5912);
	dataBufferOut(5417) <= dataBufferIn( 511) when (flag_long='1') else dataBufferIn(5995);
	dataBufferOut(5418) <= dataBufferIn(1254) when (flag_long='1') else dataBufferIn(6078);
	dataBufferOut(5419) <= dataBufferIn(1997) when (flag_long='1') else dataBufferIn(5105);
	dataBufferOut(5420) <= dataBufferIn(2740) when (flag_long='1') else dataBufferIn(5188);
	dataBufferOut(5421) <= dataBufferIn(3483) when (flag_long='1') else dataBufferIn(5271);
	dataBufferOut(5422) <= dataBufferIn(4226) when (flag_long='1') else dataBufferIn(5354);
	dataBufferOut(5423) <= dataBufferIn(4969) when (flag_long='1') else dataBufferIn(5437);
	dataBufferOut(5424) <= dataBufferIn(5712) when (flag_long='1') else dataBufferIn(5520);
	dataBufferOut(5425) <= dataBufferIn( 311) when (flag_long='1') else dataBufferIn(5603);
	dataBufferOut(5426) <= dataBufferIn(1054) when (flag_long='1') else dataBufferIn(5686);
	dataBufferOut(5427) <= dataBufferIn(1797) when (flag_long='1') else dataBufferIn(5769);
	dataBufferOut(5428) <= dataBufferIn(2540) when (flag_long='1') else dataBufferIn(5852);
	dataBufferOut(5429) <= dataBufferIn(3283) when (flag_long='1') else dataBufferIn(5935);
	dataBufferOut(5430) <= dataBufferIn(4026) when (flag_long='1') else dataBufferIn(6018);
	dataBufferOut(5431) <= dataBufferIn(4769) when (flag_long='1') else dataBufferIn(6101);
	dataBufferOut(5432) <= dataBufferIn(5512) when (flag_long='1') else dataBufferIn(5128);
	dataBufferOut(5433) <= dataBufferIn( 111) when (flag_long='1') else dataBufferIn(5211);
	dataBufferOut(5434) <= dataBufferIn( 854) when (flag_long='1') else dataBufferIn(5294);
	dataBufferOut(5435) <= dataBufferIn(1597) when (flag_long='1') else dataBufferIn(5377);
	dataBufferOut(5436) <= dataBufferIn(2340) when (flag_long='1') else dataBufferIn(5460);
	dataBufferOut(5437) <= dataBufferIn(3083) when (flag_long='1') else dataBufferIn(5543);
	dataBufferOut(5438) <= dataBufferIn(3826) when (flag_long='1') else dataBufferIn(5626);
	dataBufferOut(5439) <= dataBufferIn(4569) when (flag_long='1') else dataBufferIn(5709);
	dataBufferOut(5440) <= dataBufferIn(5312) when (flag_long='1') else dataBufferIn(5792);
	dataBufferOut(5441) <= dataBufferIn(6055) when (flag_long='1') else dataBufferIn(5875);
	dataBufferOut(5442) <= dataBufferIn( 654) when (flag_long='1') else dataBufferIn(5958);
	dataBufferOut(5443) <= dataBufferIn(1397) when (flag_long='1') else dataBufferIn(6041);
	dataBufferOut(5444) <= dataBufferIn(2140) when (flag_long='1') else dataBufferIn(6124);
	dataBufferOut(5445) <= dataBufferIn(2883) when (flag_long='1') else dataBufferIn(5151);
	dataBufferOut(5446) <= dataBufferIn(3626) when (flag_long='1') else dataBufferIn(5234);
	dataBufferOut(5447) <= dataBufferIn(4369) when (flag_long='1') else dataBufferIn(5317);
	dataBufferOut(5448) <= dataBufferIn(5112) when (flag_long='1') else dataBufferIn(5400);
	dataBufferOut(5449) <= dataBufferIn(5855) when (flag_long='1') else dataBufferIn(5483);
	dataBufferOut(5450) <= dataBufferIn( 454) when (flag_long='1') else dataBufferIn(5566);
	dataBufferOut(5451) <= dataBufferIn(1197) when (flag_long='1') else dataBufferIn(5649);
	dataBufferOut(5452) <= dataBufferIn(1940) when (flag_long='1') else dataBufferIn(5732);
	dataBufferOut(5453) <= dataBufferIn(2683) when (flag_long='1') else dataBufferIn(5815);
	dataBufferOut(5454) <= dataBufferIn(3426) when (flag_long='1') else dataBufferIn(5898);
	dataBufferOut(5455) <= dataBufferIn(4169) when (flag_long='1') else dataBufferIn(5981);
	dataBufferOut(5456) <= dataBufferIn(4912) when (flag_long='1') else dataBufferIn(6064);
	dataBufferOut(5457) <= dataBufferIn(5655) when (flag_long='1') else dataBufferIn(5091);
	dataBufferOut(5458) <= dataBufferIn( 254) when (flag_long='1') else dataBufferIn(5174);
	dataBufferOut(5459) <= dataBufferIn( 997) when (flag_long='1') else dataBufferIn(5257);
	dataBufferOut(5460) <= dataBufferIn(1740) when (flag_long='1') else dataBufferIn(5340);
	dataBufferOut(5461) <= dataBufferIn(2483) when (flag_long='1') else dataBufferIn(5423);
	dataBufferOut(5462) <= dataBufferIn(3226) when (flag_long='1') else dataBufferIn(5506);
	dataBufferOut(5463) <= dataBufferIn(3969) when (flag_long='1') else dataBufferIn(5589);
	dataBufferOut(5464) <= dataBufferIn(4712) when (flag_long='1') else dataBufferIn(5672);
	dataBufferOut(5465) <= dataBufferIn(5455) when (flag_long='1') else dataBufferIn(5755);
	dataBufferOut(5466) <= dataBufferIn(  54) when (flag_long='1') else dataBufferIn(5838);
	dataBufferOut(5467) <= dataBufferIn( 797) when (flag_long='1') else dataBufferIn(5921);
	dataBufferOut(5468) <= dataBufferIn(1540) when (flag_long='1') else dataBufferIn(6004);
	dataBufferOut(5469) <= dataBufferIn(2283) when (flag_long='1') else dataBufferIn(6087);
	dataBufferOut(5470) <= dataBufferIn(3026) when (flag_long='1') else dataBufferIn(5114);
	dataBufferOut(5471) <= dataBufferIn(3769) when (flag_long='1') else dataBufferIn(5197);
	dataBufferOut(5472) <= dataBufferIn(4512) when (flag_long='1') else dataBufferIn(5280);
	dataBufferOut(5473) <= dataBufferIn(5255) when (flag_long='1') else dataBufferIn(5363);
	dataBufferOut(5474) <= dataBufferIn(5998) when (flag_long='1') else dataBufferIn(5446);
	dataBufferOut(5475) <= dataBufferIn( 597) when (flag_long='1') else dataBufferIn(5529);
	dataBufferOut(5476) <= dataBufferIn(1340) when (flag_long='1') else dataBufferIn(5612);
	dataBufferOut(5477) <= dataBufferIn(2083) when (flag_long='1') else dataBufferIn(5695);
	dataBufferOut(5478) <= dataBufferIn(2826) when (flag_long='1') else dataBufferIn(5778);
	dataBufferOut(5479) <= dataBufferIn(3569) when (flag_long='1') else dataBufferIn(5861);
	dataBufferOut(5480) <= dataBufferIn(4312) when (flag_long='1') else dataBufferIn(5944);
	dataBufferOut(5481) <= dataBufferIn(5055) when (flag_long='1') else dataBufferIn(6027);
	dataBufferOut(5482) <= dataBufferIn(5798) when (flag_long='1') else dataBufferIn(6110);
	dataBufferOut(5483) <= dataBufferIn( 397) when (flag_long='1') else dataBufferIn(5137);
	dataBufferOut(5484) <= dataBufferIn(1140) when (flag_long='1') else dataBufferIn(5220);
	dataBufferOut(5485) <= dataBufferIn(1883) when (flag_long='1') else dataBufferIn(5303);
	dataBufferOut(5486) <= dataBufferIn(2626) when (flag_long='1') else dataBufferIn(5386);
	dataBufferOut(5487) <= dataBufferIn(3369) when (flag_long='1') else dataBufferIn(5469);
	dataBufferOut(5488) <= dataBufferIn(4112) when (flag_long='1') else dataBufferIn(5552);
	dataBufferOut(5489) <= dataBufferIn(4855) when (flag_long='1') else dataBufferIn(5635);
	dataBufferOut(5490) <= dataBufferIn(5598) when (flag_long='1') else dataBufferIn(5718);
	dataBufferOut(5491) <= dataBufferIn( 197) when (flag_long='1') else dataBufferIn(5801);
	dataBufferOut(5492) <= dataBufferIn( 940) when (flag_long='1') else dataBufferIn(5884);
	dataBufferOut(5493) <= dataBufferIn(1683) when (flag_long='1') else dataBufferIn(5967);
	dataBufferOut(5494) <= dataBufferIn(2426) when (flag_long='1') else dataBufferIn(6050);
	dataBufferOut(5495) <= dataBufferIn(3169) when (flag_long='1') else dataBufferIn(6133);
	dataBufferOut(5496) <= dataBufferIn(3912) when (flag_long='1') else dataBufferIn(5160);
	dataBufferOut(5497) <= dataBufferIn(4655) when (flag_long='1') else dataBufferIn(5243);
	dataBufferOut(5498) <= dataBufferIn(5398) when (flag_long='1') else dataBufferIn(5326);
	dataBufferOut(5499) <= dataBufferIn(6141) when (flag_long='1') else dataBufferIn(5409);
	dataBufferOut(5500) <= dataBufferIn( 740) when (flag_long='1') else dataBufferIn(5492);
	dataBufferOut(5501) <= dataBufferIn(1483) when (flag_long='1') else dataBufferIn(5575);
	dataBufferOut(5502) <= dataBufferIn(2226) when (flag_long='1') else dataBufferIn(5658);
	dataBufferOut(5503) <= dataBufferIn(2969) when (flag_long='1') else dataBufferIn(5741);
	dataBufferOut(5504) <= dataBufferIn(3712) when (flag_long='1') else dataBufferIn(5824);
	dataBufferOut(5505) <= dataBufferIn(4455) when (flag_long='1') else dataBufferIn(5907);
	dataBufferOut(5506) <= dataBufferIn(5198) when (flag_long='1') else dataBufferIn(5990);
	dataBufferOut(5507) <= dataBufferIn(5941) when (flag_long='1') else dataBufferIn(6073);
	dataBufferOut(5508) <= dataBufferIn( 540) when (flag_long='1') else dataBufferIn(5100);
	dataBufferOut(5509) <= dataBufferIn(1283) when (flag_long='1') else dataBufferIn(5183);
	dataBufferOut(5510) <= dataBufferIn(2026) when (flag_long='1') else dataBufferIn(5266);
	dataBufferOut(5511) <= dataBufferIn(2769) when (flag_long='1') else dataBufferIn(5349);
	dataBufferOut(5512) <= dataBufferIn(3512) when (flag_long='1') else dataBufferIn(5432);
	dataBufferOut(5513) <= dataBufferIn(4255) when (flag_long='1') else dataBufferIn(5515);
	dataBufferOut(5514) <= dataBufferIn(4998) when (flag_long='1') else dataBufferIn(5598);
	dataBufferOut(5515) <= dataBufferIn(5741) when (flag_long='1') else dataBufferIn(5681);
	dataBufferOut(5516) <= dataBufferIn( 340) when (flag_long='1') else dataBufferIn(5764);
	dataBufferOut(5517) <= dataBufferIn(1083) when (flag_long='1') else dataBufferIn(5847);
	dataBufferOut(5518) <= dataBufferIn(1826) when (flag_long='1') else dataBufferIn(5930);
	dataBufferOut(5519) <= dataBufferIn(2569) when (flag_long='1') else dataBufferIn(6013);
	dataBufferOut(5520) <= dataBufferIn(3312) when (flag_long='1') else dataBufferIn(6096);
	dataBufferOut(5521) <= dataBufferIn(4055) when (flag_long='1') else dataBufferIn(5123);
	dataBufferOut(5522) <= dataBufferIn(4798) when (flag_long='1') else dataBufferIn(5206);
	dataBufferOut(5523) <= dataBufferIn(5541) when (flag_long='1') else dataBufferIn(5289);
	dataBufferOut(5524) <= dataBufferIn( 140) when (flag_long='1') else dataBufferIn(5372);
	dataBufferOut(5525) <= dataBufferIn( 883) when (flag_long='1') else dataBufferIn(5455);
	dataBufferOut(5526) <= dataBufferIn(1626) when (flag_long='1') else dataBufferIn(5538);
	dataBufferOut(5527) <= dataBufferIn(2369) when (flag_long='1') else dataBufferIn(5621);
	dataBufferOut(5528) <= dataBufferIn(3112) when (flag_long='1') else dataBufferIn(5704);
	dataBufferOut(5529) <= dataBufferIn(3855) when (flag_long='1') else dataBufferIn(5787);
	dataBufferOut(5530) <= dataBufferIn(4598) when (flag_long='1') else dataBufferIn(5870);
	dataBufferOut(5531) <= dataBufferIn(5341) when (flag_long='1') else dataBufferIn(5953);
	dataBufferOut(5532) <= dataBufferIn(6084) when (flag_long='1') else dataBufferIn(6036);
	dataBufferOut(5533) <= dataBufferIn( 683) when (flag_long='1') else dataBufferIn(6119);
	dataBufferOut(5534) <= dataBufferIn(1426) when (flag_long='1') else dataBufferIn(5146);
	dataBufferOut(5535) <= dataBufferIn(2169) when (flag_long='1') else dataBufferIn(5229);
	dataBufferOut(5536) <= dataBufferIn(2912) when (flag_long='1') else dataBufferIn(5312);
	dataBufferOut(5537) <= dataBufferIn(3655) when (flag_long='1') else dataBufferIn(5395);
	dataBufferOut(5538) <= dataBufferIn(4398) when (flag_long='1') else dataBufferIn(5478);
	dataBufferOut(5539) <= dataBufferIn(5141) when (flag_long='1') else dataBufferIn(5561);
	dataBufferOut(5540) <= dataBufferIn(5884) when (flag_long='1') else dataBufferIn(5644);
	dataBufferOut(5541) <= dataBufferIn( 483) when (flag_long='1') else dataBufferIn(5727);
	dataBufferOut(5542) <= dataBufferIn(1226) when (flag_long='1') else dataBufferIn(5810);
	dataBufferOut(5543) <= dataBufferIn(1969) when (flag_long='1') else dataBufferIn(5893);
	dataBufferOut(5544) <= dataBufferIn(2712) when (flag_long='1') else dataBufferIn(5976);
	dataBufferOut(5545) <= dataBufferIn(3455) when (flag_long='1') else dataBufferIn(6059);
	dataBufferOut(5546) <= dataBufferIn(4198) when (flag_long='1') else dataBufferIn(6142);
	dataBufferOut(5547) <= dataBufferIn(4941) when (flag_long='1') else dataBufferIn(5169);
	dataBufferOut(5548) <= dataBufferIn(5684) when (flag_long='1') else dataBufferIn(5252);
	dataBufferOut(5549) <= dataBufferIn( 283) when (flag_long='1') else dataBufferIn(5335);
	dataBufferOut(5550) <= dataBufferIn(1026) when (flag_long='1') else dataBufferIn(5418);
	dataBufferOut(5551) <= dataBufferIn(1769) when (flag_long='1') else dataBufferIn(5501);
	dataBufferOut(5552) <= dataBufferIn(2512) when (flag_long='1') else dataBufferIn(5584);
	dataBufferOut(5553) <= dataBufferIn(3255) when (flag_long='1') else dataBufferIn(5667);
	dataBufferOut(5554) <= dataBufferIn(3998) when (flag_long='1') else dataBufferIn(5750);
	dataBufferOut(5555) <= dataBufferIn(4741) when (flag_long='1') else dataBufferIn(5833);
	dataBufferOut(5556) <= dataBufferIn(5484) when (flag_long='1') else dataBufferIn(5916);
	dataBufferOut(5557) <= dataBufferIn(  83) when (flag_long='1') else dataBufferIn(5999);
	dataBufferOut(5558) <= dataBufferIn( 826) when (flag_long='1') else dataBufferIn(6082);
	dataBufferOut(5559) <= dataBufferIn(1569) when (flag_long='1') else dataBufferIn(5109);
	dataBufferOut(5560) <= dataBufferIn(2312) when (flag_long='1') else dataBufferIn(5192);
	dataBufferOut(5561) <= dataBufferIn(3055) when (flag_long='1') else dataBufferIn(5275);
	dataBufferOut(5562) <= dataBufferIn(3798) when (flag_long='1') else dataBufferIn(5358);
	dataBufferOut(5563) <= dataBufferIn(4541) when (flag_long='1') else dataBufferIn(5441);
	dataBufferOut(5564) <= dataBufferIn(5284) when (flag_long='1') else dataBufferIn(5524);
	dataBufferOut(5565) <= dataBufferIn(6027) when (flag_long='1') else dataBufferIn(5607);
	dataBufferOut(5566) <= dataBufferIn( 626) when (flag_long='1') else dataBufferIn(5690);
	dataBufferOut(5567) <= dataBufferIn(1369) when (flag_long='1') else dataBufferIn(5773);
	dataBufferOut(5568) <= dataBufferIn(2112) when (flag_long='1') else dataBufferIn(5856);
	dataBufferOut(5569) <= dataBufferIn(2855) when (flag_long='1') else dataBufferIn(5939);
	dataBufferOut(5570) <= dataBufferIn(3598) when (flag_long='1') else dataBufferIn(6022);
	dataBufferOut(5571) <= dataBufferIn(4341) when (flag_long='1') else dataBufferIn(6105);
	dataBufferOut(5572) <= dataBufferIn(5084) when (flag_long='1') else dataBufferIn(5132);
	dataBufferOut(5573) <= dataBufferIn(5827) when (flag_long='1') else dataBufferIn(5215);
	dataBufferOut(5574) <= dataBufferIn( 426) when (flag_long='1') else dataBufferIn(5298);
	dataBufferOut(5575) <= dataBufferIn(1169) when (flag_long='1') else dataBufferIn(5381);
	dataBufferOut(5576) <= dataBufferIn(1912) when (flag_long='1') else dataBufferIn(5464);
	dataBufferOut(5577) <= dataBufferIn(2655) when (flag_long='1') else dataBufferIn(5547);
	dataBufferOut(5578) <= dataBufferIn(3398) when (flag_long='1') else dataBufferIn(5630);
	dataBufferOut(5579) <= dataBufferIn(4141) when (flag_long='1') else dataBufferIn(5713);
	dataBufferOut(5580) <= dataBufferIn(4884) when (flag_long='1') else dataBufferIn(5796);
	dataBufferOut(5581) <= dataBufferIn(5627) when (flag_long='1') else dataBufferIn(5879);
	dataBufferOut(5582) <= dataBufferIn( 226) when (flag_long='1') else dataBufferIn(5962);
	dataBufferOut(5583) <= dataBufferIn( 969) when (flag_long='1') else dataBufferIn(6045);
	dataBufferOut(5584) <= dataBufferIn(1712) when (flag_long='1') else dataBufferIn(6128);
	dataBufferOut(5585) <= dataBufferIn(2455) when (flag_long='1') else dataBufferIn(5155);
	dataBufferOut(5586) <= dataBufferIn(3198) when (flag_long='1') else dataBufferIn(5238);
	dataBufferOut(5587) <= dataBufferIn(3941) when (flag_long='1') else dataBufferIn(5321);
	dataBufferOut(5588) <= dataBufferIn(4684) when (flag_long='1') else dataBufferIn(5404);
	dataBufferOut(5589) <= dataBufferIn(5427) when (flag_long='1') else dataBufferIn(5487);
	dataBufferOut(5590) <= dataBufferIn(  26) when (flag_long='1') else dataBufferIn(5570);
	dataBufferOut(5591) <= dataBufferIn( 769) when (flag_long='1') else dataBufferIn(5653);
	dataBufferOut(5592) <= dataBufferIn(1512) when (flag_long='1') else dataBufferIn(5736);
	dataBufferOut(5593) <= dataBufferIn(2255) when (flag_long='1') else dataBufferIn(5819);
	dataBufferOut(5594) <= dataBufferIn(2998) when (flag_long='1') else dataBufferIn(5902);
	dataBufferOut(5595) <= dataBufferIn(3741) when (flag_long='1') else dataBufferIn(5985);
	dataBufferOut(5596) <= dataBufferIn(4484) when (flag_long='1') else dataBufferIn(6068);
	dataBufferOut(5597) <= dataBufferIn(5227) when (flag_long='1') else dataBufferIn(5095);
	dataBufferOut(5598) <= dataBufferIn(5970) when (flag_long='1') else dataBufferIn(5178);
	dataBufferOut(5599) <= dataBufferIn( 569) when (flag_long='1') else dataBufferIn(5261);
	dataBufferOut(5600) <= dataBufferIn(1312) when (flag_long='1') else dataBufferIn(5344);
	dataBufferOut(5601) <= dataBufferIn(2055) when (flag_long='1') else dataBufferIn(5427);
	dataBufferOut(5602) <= dataBufferIn(2798) when (flag_long='1') else dataBufferIn(5510);
	dataBufferOut(5603) <= dataBufferIn(3541) when (flag_long='1') else dataBufferIn(5593);
	dataBufferOut(5604) <= dataBufferIn(4284) when (flag_long='1') else dataBufferIn(5676);
	dataBufferOut(5605) <= dataBufferIn(5027) when (flag_long='1') else dataBufferIn(5759);
	dataBufferOut(5606) <= dataBufferIn(5770) when (flag_long='1') else dataBufferIn(5842);
	dataBufferOut(5607) <= dataBufferIn( 369) when (flag_long='1') else dataBufferIn(5925);
	dataBufferOut(5608) <= dataBufferIn(1112) when (flag_long='1') else dataBufferIn(6008);
	dataBufferOut(5609) <= dataBufferIn(1855) when (flag_long='1') else dataBufferIn(6091);
	dataBufferOut(5610) <= dataBufferIn(2598) when (flag_long='1') else dataBufferIn(5118);
	dataBufferOut(5611) <= dataBufferIn(3341) when (flag_long='1') else dataBufferIn(5201);
	dataBufferOut(5612) <= dataBufferIn(4084) when (flag_long='1') else dataBufferIn(5284);
	dataBufferOut(5613) <= dataBufferIn(4827) when (flag_long='1') else dataBufferIn(5367);
	dataBufferOut(5614) <= dataBufferIn(5570) when (flag_long='1') else dataBufferIn(5450);
	dataBufferOut(5615) <= dataBufferIn( 169) when (flag_long='1') else dataBufferIn(5533);
	dataBufferOut(5616) <= dataBufferIn( 912) when (flag_long='1') else dataBufferIn(5616);
	dataBufferOut(5617) <= dataBufferIn(1655) when (flag_long='1') else dataBufferIn(5699);
	dataBufferOut(5618) <= dataBufferIn(2398) when (flag_long='1') else dataBufferIn(5782);
	dataBufferOut(5619) <= dataBufferIn(3141) when (flag_long='1') else dataBufferIn(5865);
	dataBufferOut(5620) <= dataBufferIn(3884) when (flag_long='1') else dataBufferIn(5948);
	dataBufferOut(5621) <= dataBufferIn(4627) when (flag_long='1') else dataBufferIn(6031);
	dataBufferOut(5622) <= dataBufferIn(5370) when (flag_long='1') else dataBufferIn(6114);
	dataBufferOut(5623) <= dataBufferIn(6113) when (flag_long='1') else dataBufferIn(5141);
	dataBufferOut(5624) <= dataBufferIn( 712) when (flag_long='1') else dataBufferIn(5224);
	dataBufferOut(5625) <= dataBufferIn(1455) when (flag_long='1') else dataBufferIn(5307);
	dataBufferOut(5626) <= dataBufferIn(2198) when (flag_long='1') else dataBufferIn(5390);
	dataBufferOut(5627) <= dataBufferIn(2941) when (flag_long='1') else dataBufferIn(5473);
	dataBufferOut(5628) <= dataBufferIn(3684) when (flag_long='1') else dataBufferIn(5556);
	dataBufferOut(5629) <= dataBufferIn(4427) when (flag_long='1') else dataBufferIn(5639);
	dataBufferOut(5630) <= dataBufferIn(5170) when (flag_long='1') else dataBufferIn(5722);
	dataBufferOut(5631) <= dataBufferIn(5913) when (flag_long='1') else dataBufferIn(5805);
	dataBufferOut(5632) <= dataBufferIn( 512) when (flag_long='1') else dataBufferIn(5888);
	dataBufferOut(5633) <= dataBufferIn(1255) when (flag_long='1') else dataBufferIn(5971);
	dataBufferOut(5634) <= dataBufferIn(1998) when (flag_long='1') else dataBufferIn(6054);
	dataBufferOut(5635) <= dataBufferIn(2741) when (flag_long='1') else dataBufferIn(6137);
	dataBufferOut(5636) <= dataBufferIn(3484) when (flag_long='1') else dataBufferIn(5164);
	dataBufferOut(5637) <= dataBufferIn(4227) when (flag_long='1') else dataBufferIn(5247);
	dataBufferOut(5638) <= dataBufferIn(4970) when (flag_long='1') else dataBufferIn(5330);
	dataBufferOut(5639) <= dataBufferIn(5713) when (flag_long='1') else dataBufferIn(5413);
	dataBufferOut(5640) <= dataBufferIn( 312) when (flag_long='1') else dataBufferIn(5496);
	dataBufferOut(5641) <= dataBufferIn(1055) when (flag_long='1') else dataBufferIn(5579);
	dataBufferOut(5642) <= dataBufferIn(1798) when (flag_long='1') else dataBufferIn(5662);
	dataBufferOut(5643) <= dataBufferIn(2541) when (flag_long='1') else dataBufferIn(5745);
	dataBufferOut(5644) <= dataBufferIn(3284) when (flag_long='1') else dataBufferIn(5828);
	dataBufferOut(5645) <= dataBufferIn(4027) when (flag_long='1') else dataBufferIn(5911);
	dataBufferOut(5646) <= dataBufferIn(4770) when (flag_long='1') else dataBufferIn(5994);
	dataBufferOut(5647) <= dataBufferIn(5513) when (flag_long='1') else dataBufferIn(6077);
	dataBufferOut(5648) <= dataBufferIn( 112) when (flag_long='1') else dataBufferIn(5104);
	dataBufferOut(5649) <= dataBufferIn( 855) when (flag_long='1') else dataBufferIn(5187);
	dataBufferOut(5650) <= dataBufferIn(1598) when (flag_long='1') else dataBufferIn(5270);
	dataBufferOut(5651) <= dataBufferIn(2341) when (flag_long='1') else dataBufferIn(5353);
	dataBufferOut(5652) <= dataBufferIn(3084) when (flag_long='1') else dataBufferIn(5436);
	dataBufferOut(5653) <= dataBufferIn(3827) when (flag_long='1') else dataBufferIn(5519);
	dataBufferOut(5654) <= dataBufferIn(4570) when (flag_long='1') else dataBufferIn(5602);
	dataBufferOut(5655) <= dataBufferIn(5313) when (flag_long='1') else dataBufferIn(5685);
	dataBufferOut(5656) <= dataBufferIn(6056) when (flag_long='1') else dataBufferIn(5768);
	dataBufferOut(5657) <= dataBufferIn( 655) when (flag_long='1') else dataBufferIn(5851);
	dataBufferOut(5658) <= dataBufferIn(1398) when (flag_long='1') else dataBufferIn(5934);
	dataBufferOut(5659) <= dataBufferIn(2141) when (flag_long='1') else dataBufferIn(6017);
	dataBufferOut(5660) <= dataBufferIn(2884) when (flag_long='1') else dataBufferIn(6100);
	dataBufferOut(5661) <= dataBufferIn(3627) when (flag_long='1') else dataBufferIn(5127);
	dataBufferOut(5662) <= dataBufferIn(4370) when (flag_long='1') else dataBufferIn(5210);
	dataBufferOut(5663) <= dataBufferIn(5113) when (flag_long='1') else dataBufferIn(5293);
	dataBufferOut(5664) <= dataBufferIn(5856) when (flag_long='1') else dataBufferIn(5376);
	dataBufferOut(5665) <= dataBufferIn( 455) when (flag_long='1') else dataBufferIn(5459);
	dataBufferOut(5666) <= dataBufferIn(1198) when (flag_long='1') else dataBufferIn(5542);
	dataBufferOut(5667) <= dataBufferIn(1941) when (flag_long='1') else dataBufferIn(5625);
	dataBufferOut(5668) <= dataBufferIn(2684) when (flag_long='1') else dataBufferIn(5708);
	dataBufferOut(5669) <= dataBufferIn(3427) when (flag_long='1') else dataBufferIn(5791);
	dataBufferOut(5670) <= dataBufferIn(4170) when (flag_long='1') else dataBufferIn(5874);
	dataBufferOut(5671) <= dataBufferIn(4913) when (flag_long='1') else dataBufferIn(5957);
	dataBufferOut(5672) <= dataBufferIn(5656) when (flag_long='1') else dataBufferIn(6040);
	dataBufferOut(5673) <= dataBufferIn( 255) when (flag_long='1') else dataBufferIn(6123);
	dataBufferOut(5674) <= dataBufferIn( 998) when (flag_long='1') else dataBufferIn(5150);
	dataBufferOut(5675) <= dataBufferIn(1741) when (flag_long='1') else dataBufferIn(5233);
	dataBufferOut(5676) <= dataBufferIn(2484) when (flag_long='1') else dataBufferIn(5316);
	dataBufferOut(5677) <= dataBufferIn(3227) when (flag_long='1') else dataBufferIn(5399);
	dataBufferOut(5678) <= dataBufferIn(3970) when (flag_long='1') else dataBufferIn(5482);
	dataBufferOut(5679) <= dataBufferIn(4713) when (flag_long='1') else dataBufferIn(5565);
	dataBufferOut(5680) <= dataBufferIn(5456) when (flag_long='1') else dataBufferIn(5648);
	dataBufferOut(5681) <= dataBufferIn(  55) when (flag_long='1') else dataBufferIn(5731);
	dataBufferOut(5682) <= dataBufferIn( 798) when (flag_long='1') else dataBufferIn(5814);
	dataBufferOut(5683) <= dataBufferIn(1541) when (flag_long='1') else dataBufferIn(5897);
	dataBufferOut(5684) <= dataBufferIn(2284) when (flag_long='1') else dataBufferIn(5980);
	dataBufferOut(5685) <= dataBufferIn(3027) when (flag_long='1') else dataBufferIn(6063);
	dataBufferOut(5686) <= dataBufferIn(3770) when (flag_long='1') else dataBufferIn(5090);
	dataBufferOut(5687) <= dataBufferIn(4513) when (flag_long='1') else dataBufferIn(5173);
	dataBufferOut(5688) <= dataBufferIn(5256) when (flag_long='1') else dataBufferIn(5256);
	dataBufferOut(5689) <= dataBufferIn(5999) when (flag_long='1') else dataBufferIn(5339);
	dataBufferOut(5690) <= dataBufferIn( 598) when (flag_long='1') else dataBufferIn(5422);
	dataBufferOut(5691) <= dataBufferIn(1341) when (flag_long='1') else dataBufferIn(5505);
	dataBufferOut(5692) <= dataBufferIn(2084) when (flag_long='1') else dataBufferIn(5588);
	dataBufferOut(5693) <= dataBufferIn(2827) when (flag_long='1') else dataBufferIn(5671);
	dataBufferOut(5694) <= dataBufferIn(3570) when (flag_long='1') else dataBufferIn(5754);
	dataBufferOut(5695) <= dataBufferIn(4313) when (flag_long='1') else dataBufferIn(5837);
	dataBufferOut(5696) <= dataBufferIn(5056) when (flag_long='1') else dataBufferIn(5920);
	dataBufferOut(5697) <= dataBufferIn(5799) when (flag_long='1') else dataBufferIn(6003);
	dataBufferOut(5698) <= dataBufferIn( 398) when (flag_long='1') else dataBufferIn(6086);
	dataBufferOut(5699) <= dataBufferIn(1141) when (flag_long='1') else dataBufferIn(5113);
	dataBufferOut(5700) <= dataBufferIn(1884) when (flag_long='1') else dataBufferIn(5196);
	dataBufferOut(5701) <= dataBufferIn(2627) when (flag_long='1') else dataBufferIn(5279);
	dataBufferOut(5702) <= dataBufferIn(3370) when (flag_long='1') else dataBufferIn(5362);
	dataBufferOut(5703) <= dataBufferIn(4113) when (flag_long='1') else dataBufferIn(5445);
	dataBufferOut(5704) <= dataBufferIn(4856) when (flag_long='1') else dataBufferIn(5528);
	dataBufferOut(5705) <= dataBufferIn(5599) when (flag_long='1') else dataBufferIn(5611);
	dataBufferOut(5706) <= dataBufferIn( 198) when (flag_long='1') else dataBufferIn(5694);
	dataBufferOut(5707) <= dataBufferIn( 941) when (flag_long='1') else dataBufferIn(5777);
	dataBufferOut(5708) <= dataBufferIn(1684) when (flag_long='1') else dataBufferIn(5860);
	dataBufferOut(5709) <= dataBufferIn(2427) when (flag_long='1') else dataBufferIn(5943);
	dataBufferOut(5710) <= dataBufferIn(3170) when (flag_long='1') else dataBufferIn(6026);
	dataBufferOut(5711) <= dataBufferIn(3913) when (flag_long='1') else dataBufferIn(6109);
	dataBufferOut(5712) <= dataBufferIn(4656) when (flag_long='1') else dataBufferIn(5136);
	dataBufferOut(5713) <= dataBufferIn(5399) when (flag_long='1') else dataBufferIn(5219);
	dataBufferOut(5714) <= dataBufferIn(6142) when (flag_long='1') else dataBufferIn(5302);
	dataBufferOut(5715) <= dataBufferIn( 741) when (flag_long='1') else dataBufferIn(5385);
	dataBufferOut(5716) <= dataBufferIn(1484) when (flag_long='1') else dataBufferIn(5468);
	dataBufferOut(5717) <= dataBufferIn(2227) when (flag_long='1') else dataBufferIn(5551);
	dataBufferOut(5718) <= dataBufferIn(2970) when (flag_long='1') else dataBufferIn(5634);
	dataBufferOut(5719) <= dataBufferIn(3713) when (flag_long='1') else dataBufferIn(5717);
	dataBufferOut(5720) <= dataBufferIn(4456) when (flag_long='1') else dataBufferIn(5800);
	dataBufferOut(5721) <= dataBufferIn(5199) when (flag_long='1') else dataBufferIn(5883);
	dataBufferOut(5722) <= dataBufferIn(5942) when (flag_long='1') else dataBufferIn(5966);
	dataBufferOut(5723) <= dataBufferIn( 541) when (flag_long='1') else dataBufferIn(6049);
	dataBufferOut(5724) <= dataBufferIn(1284) when (flag_long='1') else dataBufferIn(6132);
	dataBufferOut(5725) <= dataBufferIn(2027) when (flag_long='1') else dataBufferIn(5159);
	dataBufferOut(5726) <= dataBufferIn(2770) when (flag_long='1') else dataBufferIn(5242);
	dataBufferOut(5727) <= dataBufferIn(3513) when (flag_long='1') else dataBufferIn(5325);
	dataBufferOut(5728) <= dataBufferIn(4256) when (flag_long='1') else dataBufferIn(5408);
	dataBufferOut(5729) <= dataBufferIn(4999) when (flag_long='1') else dataBufferIn(5491);
	dataBufferOut(5730) <= dataBufferIn(5742) when (flag_long='1') else dataBufferIn(5574);
	dataBufferOut(5731) <= dataBufferIn( 341) when (flag_long='1') else dataBufferIn(5657);
	dataBufferOut(5732) <= dataBufferIn(1084) when (flag_long='1') else dataBufferIn(5740);
	dataBufferOut(5733) <= dataBufferIn(1827) when (flag_long='1') else dataBufferIn(5823);
	dataBufferOut(5734) <= dataBufferIn(2570) when (flag_long='1') else dataBufferIn(5906);
	dataBufferOut(5735) <= dataBufferIn(3313) when (flag_long='1') else dataBufferIn(5989);
	dataBufferOut(5736) <= dataBufferIn(4056) when (flag_long='1') else dataBufferIn(6072);
	dataBufferOut(5737) <= dataBufferIn(4799) when (flag_long='1') else dataBufferIn(5099);
	dataBufferOut(5738) <= dataBufferIn(5542) when (flag_long='1') else dataBufferIn(5182);
	dataBufferOut(5739) <= dataBufferIn( 141) when (flag_long='1') else dataBufferIn(5265);
	dataBufferOut(5740) <= dataBufferIn( 884) when (flag_long='1') else dataBufferIn(5348);
	dataBufferOut(5741) <= dataBufferIn(1627) when (flag_long='1') else dataBufferIn(5431);
	dataBufferOut(5742) <= dataBufferIn(2370) when (flag_long='1') else dataBufferIn(5514);
	dataBufferOut(5743) <= dataBufferIn(3113) when (flag_long='1') else dataBufferIn(5597);
	dataBufferOut(5744) <= dataBufferIn(3856) when (flag_long='1') else dataBufferIn(5680);
	dataBufferOut(5745) <= dataBufferIn(4599) when (flag_long='1') else dataBufferIn(5763);
	dataBufferOut(5746) <= dataBufferIn(5342) when (flag_long='1') else dataBufferIn(5846);
	dataBufferOut(5747) <= dataBufferIn(6085) when (flag_long='1') else dataBufferIn(5929);
	dataBufferOut(5748) <= dataBufferIn( 684) when (flag_long='1') else dataBufferIn(6012);
	dataBufferOut(5749) <= dataBufferIn(1427) when (flag_long='1') else dataBufferIn(6095);
	dataBufferOut(5750) <= dataBufferIn(2170) when (flag_long='1') else dataBufferIn(5122);
	dataBufferOut(5751) <= dataBufferIn(2913) when (flag_long='1') else dataBufferIn(5205);
	dataBufferOut(5752) <= dataBufferIn(3656) when (flag_long='1') else dataBufferIn(5288);
	dataBufferOut(5753) <= dataBufferIn(4399) when (flag_long='1') else dataBufferIn(5371);
	dataBufferOut(5754) <= dataBufferIn(5142) when (flag_long='1') else dataBufferIn(5454);
	dataBufferOut(5755) <= dataBufferIn(5885) when (flag_long='1') else dataBufferIn(5537);
	dataBufferOut(5756) <= dataBufferIn( 484) when (flag_long='1') else dataBufferIn(5620);
	dataBufferOut(5757) <= dataBufferIn(1227) when (flag_long='1') else dataBufferIn(5703);
	dataBufferOut(5758) <= dataBufferIn(1970) when (flag_long='1') else dataBufferIn(5786);
	dataBufferOut(5759) <= dataBufferIn(2713) when (flag_long='1') else dataBufferIn(5869);
	dataBufferOut(5760) <= dataBufferIn(3456) when (flag_long='1') else dataBufferIn(5952);
	dataBufferOut(5761) <= dataBufferIn(4199) when (flag_long='1') else dataBufferIn(6035);
	dataBufferOut(5762) <= dataBufferIn(4942) when (flag_long='1') else dataBufferIn(6118);
	dataBufferOut(5763) <= dataBufferIn(5685) when (flag_long='1') else dataBufferIn(5145);
	dataBufferOut(5764) <= dataBufferIn( 284) when (flag_long='1') else dataBufferIn(5228);
	dataBufferOut(5765) <= dataBufferIn(1027) when (flag_long='1') else dataBufferIn(5311);
	dataBufferOut(5766) <= dataBufferIn(1770) when (flag_long='1') else dataBufferIn(5394);
	dataBufferOut(5767) <= dataBufferIn(2513) when (flag_long='1') else dataBufferIn(5477);
	dataBufferOut(5768) <= dataBufferIn(3256) when (flag_long='1') else dataBufferIn(5560);
	dataBufferOut(5769) <= dataBufferIn(3999) when (flag_long='1') else dataBufferIn(5643);
	dataBufferOut(5770) <= dataBufferIn(4742) when (flag_long='1') else dataBufferIn(5726);
	dataBufferOut(5771) <= dataBufferIn(5485) when (flag_long='1') else dataBufferIn(5809);
	dataBufferOut(5772) <= dataBufferIn(  84) when (flag_long='1') else dataBufferIn(5892);
	dataBufferOut(5773) <= dataBufferIn( 827) when (flag_long='1') else dataBufferIn(5975);
	dataBufferOut(5774) <= dataBufferIn(1570) when (flag_long='1') else dataBufferIn(6058);
	dataBufferOut(5775) <= dataBufferIn(2313) when (flag_long='1') else dataBufferIn(6141);
	dataBufferOut(5776) <= dataBufferIn(3056) when (flag_long='1') else dataBufferIn(5168);
	dataBufferOut(5777) <= dataBufferIn(3799) when (flag_long='1') else dataBufferIn(5251);
	dataBufferOut(5778) <= dataBufferIn(4542) when (flag_long='1') else dataBufferIn(5334);
	dataBufferOut(5779) <= dataBufferIn(5285) when (flag_long='1') else dataBufferIn(5417);
	dataBufferOut(5780) <= dataBufferIn(6028) when (flag_long='1') else dataBufferIn(5500);
	dataBufferOut(5781) <= dataBufferIn( 627) when (flag_long='1') else dataBufferIn(5583);
	dataBufferOut(5782) <= dataBufferIn(1370) when (flag_long='1') else dataBufferIn(5666);
	dataBufferOut(5783) <= dataBufferIn(2113) when (flag_long='1') else dataBufferIn(5749);
	dataBufferOut(5784) <= dataBufferIn(2856) when (flag_long='1') else dataBufferIn(5832);
	dataBufferOut(5785) <= dataBufferIn(3599) when (flag_long='1') else dataBufferIn(5915);
	dataBufferOut(5786) <= dataBufferIn(4342) when (flag_long='1') else dataBufferIn(5998);
	dataBufferOut(5787) <= dataBufferIn(5085) when (flag_long='1') else dataBufferIn(6081);
	dataBufferOut(5788) <= dataBufferIn(5828) when (flag_long='1') else dataBufferIn(5108);
	dataBufferOut(5789) <= dataBufferIn( 427) when (flag_long='1') else dataBufferIn(5191);
	dataBufferOut(5790) <= dataBufferIn(1170) when (flag_long='1') else dataBufferIn(5274);
	dataBufferOut(5791) <= dataBufferIn(1913) when (flag_long='1') else dataBufferIn(5357);
	dataBufferOut(5792) <= dataBufferIn(2656) when (flag_long='1') else dataBufferIn(5440);
	dataBufferOut(5793) <= dataBufferIn(3399) when (flag_long='1') else dataBufferIn(5523);
	dataBufferOut(5794) <= dataBufferIn(4142) when (flag_long='1') else dataBufferIn(5606);
	dataBufferOut(5795) <= dataBufferIn(4885) when (flag_long='1') else dataBufferIn(5689);
	dataBufferOut(5796) <= dataBufferIn(5628) when (flag_long='1') else dataBufferIn(5772);
	dataBufferOut(5797) <= dataBufferIn( 227) when (flag_long='1') else dataBufferIn(5855);
	dataBufferOut(5798) <= dataBufferIn( 970) when (flag_long='1') else dataBufferIn(5938);
	dataBufferOut(5799) <= dataBufferIn(1713) when (flag_long='1') else dataBufferIn(6021);
	dataBufferOut(5800) <= dataBufferIn(2456) when (flag_long='1') else dataBufferIn(6104);
	dataBufferOut(5801) <= dataBufferIn(3199) when (flag_long='1') else dataBufferIn(5131);
	dataBufferOut(5802) <= dataBufferIn(3942) when (flag_long='1') else dataBufferIn(5214);
	dataBufferOut(5803) <= dataBufferIn(4685) when (flag_long='1') else dataBufferIn(5297);
	dataBufferOut(5804) <= dataBufferIn(5428) when (flag_long='1') else dataBufferIn(5380);
	dataBufferOut(5805) <= dataBufferIn(  27) when (flag_long='1') else dataBufferIn(5463);
	dataBufferOut(5806) <= dataBufferIn( 770) when (flag_long='1') else dataBufferIn(5546);
	dataBufferOut(5807) <= dataBufferIn(1513) when (flag_long='1') else dataBufferIn(5629);
	dataBufferOut(5808) <= dataBufferIn(2256) when (flag_long='1') else dataBufferIn(5712);
	dataBufferOut(5809) <= dataBufferIn(2999) when (flag_long='1') else dataBufferIn(5795);
	dataBufferOut(5810) <= dataBufferIn(3742) when (flag_long='1') else dataBufferIn(5878);
	dataBufferOut(5811) <= dataBufferIn(4485) when (flag_long='1') else dataBufferIn(5961);
	dataBufferOut(5812) <= dataBufferIn(5228) when (flag_long='1') else dataBufferIn(6044);
	dataBufferOut(5813) <= dataBufferIn(5971) when (flag_long='1') else dataBufferIn(6127);
	dataBufferOut(5814) <= dataBufferIn( 570) when (flag_long='1') else dataBufferIn(5154);
	dataBufferOut(5815) <= dataBufferIn(1313) when (flag_long='1') else dataBufferIn(5237);
	dataBufferOut(5816) <= dataBufferIn(2056) when (flag_long='1') else dataBufferIn(5320);
	dataBufferOut(5817) <= dataBufferIn(2799) when (flag_long='1') else dataBufferIn(5403);
	dataBufferOut(5818) <= dataBufferIn(3542) when (flag_long='1') else dataBufferIn(5486);
	dataBufferOut(5819) <= dataBufferIn(4285) when (flag_long='1') else dataBufferIn(5569);
	dataBufferOut(5820) <= dataBufferIn(5028) when (flag_long='1') else dataBufferIn(5652);
	dataBufferOut(5821) <= dataBufferIn(5771) when (flag_long='1') else dataBufferIn(5735);
	dataBufferOut(5822) <= dataBufferIn( 370) when (flag_long='1') else dataBufferIn(5818);
	dataBufferOut(5823) <= dataBufferIn(1113) when (flag_long='1') else dataBufferIn(5901);
	dataBufferOut(5824) <= dataBufferIn(1856) when (flag_long='1') else dataBufferIn(5984);
	dataBufferOut(5825) <= dataBufferIn(2599) when (flag_long='1') else dataBufferIn(6067);
	dataBufferOut(5826) <= dataBufferIn(3342) when (flag_long='1') else dataBufferIn(5094);
	dataBufferOut(5827) <= dataBufferIn(4085) when (flag_long='1') else dataBufferIn(5177);
	dataBufferOut(5828) <= dataBufferIn(4828) when (flag_long='1') else dataBufferIn(5260);
	dataBufferOut(5829) <= dataBufferIn(5571) when (flag_long='1') else dataBufferIn(5343);
	dataBufferOut(5830) <= dataBufferIn( 170) when (flag_long='1') else dataBufferIn(5426);
	dataBufferOut(5831) <= dataBufferIn( 913) when (flag_long='1') else dataBufferIn(5509);
	dataBufferOut(5832) <= dataBufferIn(1656) when (flag_long='1') else dataBufferIn(5592);
	dataBufferOut(5833) <= dataBufferIn(2399) when (flag_long='1') else dataBufferIn(5675);
	dataBufferOut(5834) <= dataBufferIn(3142) when (flag_long='1') else dataBufferIn(5758);
	dataBufferOut(5835) <= dataBufferIn(3885) when (flag_long='1') else dataBufferIn(5841);
	dataBufferOut(5836) <= dataBufferIn(4628) when (flag_long='1') else dataBufferIn(5924);
	dataBufferOut(5837) <= dataBufferIn(5371) when (flag_long='1') else dataBufferIn(6007);
	dataBufferOut(5838) <= dataBufferIn(6114) when (flag_long='1') else dataBufferIn(6090);
	dataBufferOut(5839) <= dataBufferIn( 713) when (flag_long='1') else dataBufferIn(5117);
	dataBufferOut(5840) <= dataBufferIn(1456) when (flag_long='1') else dataBufferIn(5200);
	dataBufferOut(5841) <= dataBufferIn(2199) when (flag_long='1') else dataBufferIn(5283);
	dataBufferOut(5842) <= dataBufferIn(2942) when (flag_long='1') else dataBufferIn(5366);
	dataBufferOut(5843) <= dataBufferIn(3685) when (flag_long='1') else dataBufferIn(5449);
	dataBufferOut(5844) <= dataBufferIn(4428) when (flag_long='1') else dataBufferIn(5532);
	dataBufferOut(5845) <= dataBufferIn(5171) when (flag_long='1') else dataBufferIn(5615);
	dataBufferOut(5846) <= dataBufferIn(5914) when (flag_long='1') else dataBufferIn(5698);
	dataBufferOut(5847) <= dataBufferIn( 513) when (flag_long='1') else dataBufferIn(5781);
	dataBufferOut(5848) <= dataBufferIn(1256) when (flag_long='1') else dataBufferIn(5864);
	dataBufferOut(5849) <= dataBufferIn(1999) when (flag_long='1') else dataBufferIn(5947);
	dataBufferOut(5850) <= dataBufferIn(2742) when (flag_long='1') else dataBufferIn(6030);
	dataBufferOut(5851) <= dataBufferIn(3485) when (flag_long='1') else dataBufferIn(6113);
	dataBufferOut(5852) <= dataBufferIn(4228) when (flag_long='1') else dataBufferIn(5140);
	dataBufferOut(5853) <= dataBufferIn(4971) when (flag_long='1') else dataBufferIn(5223);
	dataBufferOut(5854) <= dataBufferIn(5714) when (flag_long='1') else dataBufferIn(5306);
	dataBufferOut(5855) <= dataBufferIn( 313) when (flag_long='1') else dataBufferIn(5389);
	dataBufferOut(5856) <= dataBufferIn(1056) when (flag_long='1') else dataBufferIn(5472);
	dataBufferOut(5857) <= dataBufferIn(1799) when (flag_long='1') else dataBufferIn(5555);
	dataBufferOut(5858) <= dataBufferIn(2542) when (flag_long='1') else dataBufferIn(5638);
	dataBufferOut(5859) <= dataBufferIn(3285) when (flag_long='1') else dataBufferIn(5721);
	dataBufferOut(5860) <= dataBufferIn(4028) when (flag_long='1') else dataBufferIn(5804);
	dataBufferOut(5861) <= dataBufferIn(4771) when (flag_long='1') else dataBufferIn(5887);
	dataBufferOut(5862) <= dataBufferIn(5514) when (flag_long='1') else dataBufferIn(5970);
	dataBufferOut(5863) <= dataBufferIn( 113) when (flag_long='1') else dataBufferIn(6053);
	dataBufferOut(5864) <= dataBufferIn( 856) when (flag_long='1') else dataBufferIn(6136);
	dataBufferOut(5865) <= dataBufferIn(1599) when (flag_long='1') else dataBufferIn(5163);
	dataBufferOut(5866) <= dataBufferIn(2342) when (flag_long='1') else dataBufferIn(5246);
	dataBufferOut(5867) <= dataBufferIn(3085) when (flag_long='1') else dataBufferIn(5329);
	dataBufferOut(5868) <= dataBufferIn(3828) when (flag_long='1') else dataBufferIn(5412);
	dataBufferOut(5869) <= dataBufferIn(4571) when (flag_long='1') else dataBufferIn(5495);
	dataBufferOut(5870) <= dataBufferIn(5314) when (flag_long='1') else dataBufferIn(5578);
	dataBufferOut(5871) <= dataBufferIn(6057) when (flag_long='1') else dataBufferIn(5661);
	dataBufferOut(5872) <= dataBufferIn( 656) when (flag_long='1') else dataBufferIn(5744);
	dataBufferOut(5873) <= dataBufferIn(1399) when (flag_long='1') else dataBufferIn(5827);
	dataBufferOut(5874) <= dataBufferIn(2142) when (flag_long='1') else dataBufferIn(5910);
	dataBufferOut(5875) <= dataBufferIn(2885) when (flag_long='1') else dataBufferIn(5993);
	dataBufferOut(5876) <= dataBufferIn(3628) when (flag_long='1') else dataBufferIn(6076);
	dataBufferOut(5877) <= dataBufferIn(4371) when (flag_long='1') else dataBufferIn(5103);
	dataBufferOut(5878) <= dataBufferIn(5114) when (flag_long='1') else dataBufferIn(5186);
	dataBufferOut(5879) <= dataBufferIn(5857) when (flag_long='1') else dataBufferIn(5269);
	dataBufferOut(5880) <= dataBufferIn( 456) when (flag_long='1') else dataBufferIn(5352);
	dataBufferOut(5881) <= dataBufferIn(1199) when (flag_long='1') else dataBufferIn(5435);
	dataBufferOut(5882) <= dataBufferIn(1942) when (flag_long='1') else dataBufferIn(5518);
	dataBufferOut(5883) <= dataBufferIn(2685) when (flag_long='1') else dataBufferIn(5601);
	dataBufferOut(5884) <= dataBufferIn(3428) when (flag_long='1') else dataBufferIn(5684);
	dataBufferOut(5885) <= dataBufferIn(4171) when (flag_long='1') else dataBufferIn(5767);
	dataBufferOut(5886) <= dataBufferIn(4914) when (flag_long='1') else dataBufferIn(5850);
	dataBufferOut(5887) <= dataBufferIn(5657) when (flag_long='1') else dataBufferIn(5933);
	dataBufferOut(5888) <= dataBufferIn( 256) when (flag_long='1') else dataBufferIn(6016);
	dataBufferOut(5889) <= dataBufferIn( 999) when (flag_long='1') else dataBufferIn(6099);
	dataBufferOut(5890) <= dataBufferIn(1742) when (flag_long='1') else dataBufferIn(5126);
	dataBufferOut(5891) <= dataBufferIn(2485) when (flag_long='1') else dataBufferIn(5209);
	dataBufferOut(5892) <= dataBufferIn(3228) when (flag_long='1') else dataBufferIn(5292);
	dataBufferOut(5893) <= dataBufferIn(3971) when (flag_long='1') else dataBufferIn(5375);
	dataBufferOut(5894) <= dataBufferIn(4714) when (flag_long='1') else dataBufferIn(5458);
	dataBufferOut(5895) <= dataBufferIn(5457) when (flag_long='1') else dataBufferIn(5541);
	dataBufferOut(5896) <= dataBufferIn(  56) when (flag_long='1') else dataBufferIn(5624);
	dataBufferOut(5897) <= dataBufferIn( 799) when (flag_long='1') else dataBufferIn(5707);
	dataBufferOut(5898) <= dataBufferIn(1542) when (flag_long='1') else dataBufferIn(5790);
	dataBufferOut(5899) <= dataBufferIn(2285) when (flag_long='1') else dataBufferIn(5873);
	dataBufferOut(5900) <= dataBufferIn(3028) when (flag_long='1') else dataBufferIn(5956);
	dataBufferOut(5901) <= dataBufferIn(3771) when (flag_long='1') else dataBufferIn(6039);
	dataBufferOut(5902) <= dataBufferIn(4514) when (flag_long='1') else dataBufferIn(6122);
	dataBufferOut(5903) <= dataBufferIn(5257) when (flag_long='1') else dataBufferIn(5149);
	dataBufferOut(5904) <= dataBufferIn(6000) when (flag_long='1') else dataBufferIn(5232);
	dataBufferOut(5905) <= dataBufferIn( 599) when (flag_long='1') else dataBufferIn(5315);
	dataBufferOut(5906) <= dataBufferIn(1342) when (flag_long='1') else dataBufferIn(5398);
	dataBufferOut(5907) <= dataBufferIn(2085) when (flag_long='1') else dataBufferIn(5481);
	dataBufferOut(5908) <= dataBufferIn(2828) when (flag_long='1') else dataBufferIn(5564);
	dataBufferOut(5909) <= dataBufferIn(3571) when (flag_long='1') else dataBufferIn(5647);
	dataBufferOut(5910) <= dataBufferIn(4314) when (flag_long='1') else dataBufferIn(5730);
	dataBufferOut(5911) <= dataBufferIn(5057) when (flag_long='1') else dataBufferIn(5813);
	dataBufferOut(5912) <= dataBufferIn(5800) when (flag_long='1') else dataBufferIn(5896);
	dataBufferOut(5913) <= dataBufferIn( 399) when (flag_long='1') else dataBufferIn(5979);
	dataBufferOut(5914) <= dataBufferIn(1142) when (flag_long='1') else dataBufferIn(6062);
	dataBufferOut(5915) <= dataBufferIn(1885) when (flag_long='1') else dataBufferIn(5089);
	dataBufferOut(5916) <= dataBufferIn(2628) when (flag_long='1') else dataBufferIn(5172);
	dataBufferOut(5917) <= dataBufferIn(3371) when (flag_long='1') else dataBufferIn(5255);
	dataBufferOut(5918) <= dataBufferIn(4114) when (flag_long='1') else dataBufferIn(5338);
	dataBufferOut(5919) <= dataBufferIn(4857) when (flag_long='1') else dataBufferIn(5421);
	dataBufferOut(5920) <= dataBufferIn(5600) when (flag_long='1') else dataBufferIn(5504);
	dataBufferOut(5921) <= dataBufferIn( 199) when (flag_long='1') else dataBufferIn(5587);
	dataBufferOut(5922) <= dataBufferIn( 942) when (flag_long='1') else dataBufferIn(5670);
	dataBufferOut(5923) <= dataBufferIn(1685) when (flag_long='1') else dataBufferIn(5753);
	dataBufferOut(5924) <= dataBufferIn(2428) when (flag_long='1') else dataBufferIn(5836);
	dataBufferOut(5925) <= dataBufferIn(3171) when (flag_long='1') else dataBufferIn(5919);
	dataBufferOut(5926) <= dataBufferIn(3914) when (flag_long='1') else dataBufferIn(6002);
	dataBufferOut(5927) <= dataBufferIn(4657) when (flag_long='1') else dataBufferIn(6085);
	dataBufferOut(5928) <= dataBufferIn(5400) when (flag_long='1') else dataBufferIn(5112);
	dataBufferOut(5929) <= dataBufferIn(6143) when (flag_long='1') else dataBufferIn(5195);
	dataBufferOut(5930) <= dataBufferIn( 742) when (flag_long='1') else dataBufferIn(5278);
	dataBufferOut(5931) <= dataBufferIn(1485) when (flag_long='1') else dataBufferIn(5361);
	dataBufferOut(5932) <= dataBufferIn(2228) when (flag_long='1') else dataBufferIn(5444);
	dataBufferOut(5933) <= dataBufferIn(2971) when (flag_long='1') else dataBufferIn(5527);
	dataBufferOut(5934) <= dataBufferIn(3714) when (flag_long='1') else dataBufferIn(5610);
	dataBufferOut(5935) <= dataBufferIn(4457) when (flag_long='1') else dataBufferIn(5693);
	dataBufferOut(5936) <= dataBufferIn(5200) when (flag_long='1') else dataBufferIn(5776);
	dataBufferOut(5937) <= dataBufferIn(5943) when (flag_long='1') else dataBufferIn(5859);
	dataBufferOut(5938) <= dataBufferIn( 542) when (flag_long='1') else dataBufferIn(5942);
	dataBufferOut(5939) <= dataBufferIn(1285) when (flag_long='1') else dataBufferIn(6025);
	dataBufferOut(5940) <= dataBufferIn(2028) when (flag_long='1') else dataBufferIn(6108);
	dataBufferOut(5941) <= dataBufferIn(2771) when (flag_long='1') else dataBufferIn(5135);
	dataBufferOut(5942) <= dataBufferIn(3514) when (flag_long='1') else dataBufferIn(5218);
	dataBufferOut(5943) <= dataBufferIn(4257) when (flag_long='1') else dataBufferIn(5301);
	dataBufferOut(5944) <= dataBufferIn(5000) when (flag_long='1') else dataBufferIn(5384);
	dataBufferOut(5945) <= dataBufferIn(5743) when (flag_long='1') else dataBufferIn(5467);
	dataBufferOut(5946) <= dataBufferIn( 342) when (flag_long='1') else dataBufferIn(5550);
	dataBufferOut(5947) <= dataBufferIn(1085) when (flag_long='1') else dataBufferIn(5633);
	dataBufferOut(5948) <= dataBufferIn(1828) when (flag_long='1') else dataBufferIn(5716);
	dataBufferOut(5949) <= dataBufferIn(2571) when (flag_long='1') else dataBufferIn(5799);
	dataBufferOut(5950) <= dataBufferIn(3314) when (flag_long='1') else dataBufferIn(5882);
	dataBufferOut(5951) <= dataBufferIn(4057) when (flag_long='1') else dataBufferIn(5965);
	dataBufferOut(5952) <= dataBufferIn(4800) when (flag_long='1') else dataBufferIn(6048);
	dataBufferOut(5953) <= dataBufferIn(5543) when (flag_long='1') else dataBufferIn(6131);
	dataBufferOut(5954) <= dataBufferIn( 142) when (flag_long='1') else dataBufferIn(5158);
	dataBufferOut(5955) <= dataBufferIn( 885) when (flag_long='1') else dataBufferIn(5241);
	dataBufferOut(5956) <= dataBufferIn(1628) when (flag_long='1') else dataBufferIn(5324);
	dataBufferOut(5957) <= dataBufferIn(2371) when (flag_long='1') else dataBufferIn(5407);
	dataBufferOut(5958) <= dataBufferIn(3114) when (flag_long='1') else dataBufferIn(5490);
	dataBufferOut(5959) <= dataBufferIn(3857) when (flag_long='1') else dataBufferIn(5573);
	dataBufferOut(5960) <= dataBufferIn(4600) when (flag_long='1') else dataBufferIn(5656);
	dataBufferOut(5961) <= dataBufferIn(5343) when (flag_long='1') else dataBufferIn(5739);
	dataBufferOut(5962) <= dataBufferIn(6086) when (flag_long='1') else dataBufferIn(5822);
	dataBufferOut(5963) <= dataBufferIn( 685) when (flag_long='1') else dataBufferIn(5905);
	dataBufferOut(5964) <= dataBufferIn(1428) when (flag_long='1') else dataBufferIn(5988);
	dataBufferOut(5965) <= dataBufferIn(2171) when (flag_long='1') else dataBufferIn(6071);
	dataBufferOut(5966) <= dataBufferIn(2914) when (flag_long='1') else dataBufferIn(5098);
	dataBufferOut(5967) <= dataBufferIn(3657) when (flag_long='1') else dataBufferIn(5181);
	dataBufferOut(5968) <= dataBufferIn(4400) when (flag_long='1') else dataBufferIn(5264);
	dataBufferOut(5969) <= dataBufferIn(5143) when (flag_long='1') else dataBufferIn(5347);
	dataBufferOut(5970) <= dataBufferIn(5886) when (flag_long='1') else dataBufferIn(5430);
	dataBufferOut(5971) <= dataBufferIn( 485) when (flag_long='1') else dataBufferIn(5513);
	dataBufferOut(5972) <= dataBufferIn(1228) when (flag_long='1') else dataBufferIn(5596);
	dataBufferOut(5973) <= dataBufferIn(1971) when (flag_long='1') else dataBufferIn(5679);
	dataBufferOut(5974) <= dataBufferIn(2714) when (flag_long='1') else dataBufferIn(5762);
	dataBufferOut(5975) <= dataBufferIn(3457) when (flag_long='1') else dataBufferIn(5845);
	dataBufferOut(5976) <= dataBufferIn(4200) when (flag_long='1') else dataBufferIn(5928);
	dataBufferOut(5977) <= dataBufferIn(4943) when (flag_long='1') else dataBufferIn(6011);
	dataBufferOut(5978) <= dataBufferIn(5686) when (flag_long='1') else dataBufferIn(6094);
	dataBufferOut(5979) <= dataBufferIn( 285) when (flag_long='1') else dataBufferIn(5121);
	dataBufferOut(5980) <= dataBufferIn(1028) when (flag_long='1') else dataBufferIn(5204);
	dataBufferOut(5981) <= dataBufferIn(1771) when (flag_long='1') else dataBufferIn(5287);
	dataBufferOut(5982) <= dataBufferIn(2514) when (flag_long='1') else dataBufferIn(5370);
	dataBufferOut(5983) <= dataBufferIn(3257) when (flag_long='1') else dataBufferIn(5453);
	dataBufferOut(5984) <= dataBufferIn(4000) when (flag_long='1') else dataBufferIn(5536);
	dataBufferOut(5985) <= dataBufferIn(4743) when (flag_long='1') else dataBufferIn(5619);
	dataBufferOut(5986) <= dataBufferIn(5486) when (flag_long='1') else dataBufferIn(5702);
	dataBufferOut(5987) <= dataBufferIn(  85) when (flag_long='1') else dataBufferIn(5785);
	dataBufferOut(5988) <= dataBufferIn( 828) when (flag_long='1') else dataBufferIn(5868);
	dataBufferOut(5989) <= dataBufferIn(1571) when (flag_long='1') else dataBufferIn(5951);
	dataBufferOut(5990) <= dataBufferIn(2314) when (flag_long='1') else dataBufferIn(6034);
	dataBufferOut(5991) <= dataBufferIn(3057) when (flag_long='1') else dataBufferIn(6117);
	dataBufferOut(5992) <= dataBufferIn(3800) when (flag_long='1') else dataBufferIn(5144);
	dataBufferOut(5993) <= dataBufferIn(4543) when (flag_long='1') else dataBufferIn(5227);
	dataBufferOut(5994) <= dataBufferIn(5286) when (flag_long='1') else dataBufferIn(5310);
	dataBufferOut(5995) <= dataBufferIn(6029) when (flag_long='1') else dataBufferIn(5393);
	dataBufferOut(5996) <= dataBufferIn( 628) when (flag_long='1') else dataBufferIn(5476);
	dataBufferOut(5997) <= dataBufferIn(1371) when (flag_long='1') else dataBufferIn(5559);
	dataBufferOut(5998) <= dataBufferIn(2114) when (flag_long='1') else dataBufferIn(5642);
	dataBufferOut(5999) <= dataBufferIn(2857) when (flag_long='1') else dataBufferIn(5725);
	dataBufferOut(6000) <= dataBufferIn(3600) when (flag_long='1') else dataBufferIn(5808);
	dataBufferOut(6001) <= dataBufferIn(4343) when (flag_long='1') else dataBufferIn(5891);
	dataBufferOut(6002) <= dataBufferIn(5086) when (flag_long='1') else dataBufferIn(5974);
	dataBufferOut(6003) <= dataBufferIn(5829) when (flag_long='1') else dataBufferIn(6057);
	dataBufferOut(6004) <= dataBufferIn( 428) when (flag_long='1') else dataBufferIn(6140);
	dataBufferOut(6005) <= dataBufferIn(1171) when (flag_long='1') else dataBufferIn(5167);
	dataBufferOut(6006) <= dataBufferIn(1914) when (flag_long='1') else dataBufferIn(5250);
	dataBufferOut(6007) <= dataBufferIn(2657) when (flag_long='1') else dataBufferIn(5333);
	dataBufferOut(6008) <= dataBufferIn(3400) when (flag_long='1') else dataBufferIn(5416);
	dataBufferOut(6009) <= dataBufferIn(4143) when (flag_long='1') else dataBufferIn(5499);
	dataBufferOut(6010) <= dataBufferIn(4886) when (flag_long='1') else dataBufferIn(5582);
	dataBufferOut(6011) <= dataBufferIn(5629) when (flag_long='1') else dataBufferIn(5665);
	dataBufferOut(6012) <= dataBufferIn( 228) when (flag_long='1') else dataBufferIn(5748);
	dataBufferOut(6013) <= dataBufferIn( 971) when (flag_long='1') else dataBufferIn(5831);
	dataBufferOut(6014) <= dataBufferIn(1714) when (flag_long='1') else dataBufferIn(5914);
	dataBufferOut(6015) <= dataBufferIn(2457) when (flag_long='1') else dataBufferIn(5997);
	dataBufferOut(6016) <= dataBufferIn(3200) when (flag_long='1') else dataBufferIn(6080);
	dataBufferOut(6017) <= dataBufferIn(3943) when (flag_long='1') else dataBufferIn(5107);
	dataBufferOut(6018) <= dataBufferIn(4686) when (flag_long='1') else dataBufferIn(5190);
	dataBufferOut(6019) <= dataBufferIn(5429) when (flag_long='1') else dataBufferIn(5273);
	dataBufferOut(6020) <= dataBufferIn(  28) when (flag_long='1') else dataBufferIn(5356);
	dataBufferOut(6021) <= dataBufferIn( 771) when (flag_long='1') else dataBufferIn(5439);
	dataBufferOut(6022) <= dataBufferIn(1514) when (flag_long='1') else dataBufferIn(5522);
	dataBufferOut(6023) <= dataBufferIn(2257) when (flag_long='1') else dataBufferIn(5605);
	dataBufferOut(6024) <= dataBufferIn(3000) when (flag_long='1') else dataBufferIn(5688);
	dataBufferOut(6025) <= dataBufferIn(3743) when (flag_long='1') else dataBufferIn(5771);
	dataBufferOut(6026) <= dataBufferIn(4486) when (flag_long='1') else dataBufferIn(5854);
	dataBufferOut(6027) <= dataBufferIn(5229) when (flag_long='1') else dataBufferIn(5937);
	dataBufferOut(6028) <= dataBufferIn(5972) when (flag_long='1') else dataBufferIn(6020);
	dataBufferOut(6029) <= dataBufferIn( 571) when (flag_long='1') else dataBufferIn(6103);
	dataBufferOut(6030) <= dataBufferIn(1314) when (flag_long='1') else dataBufferIn(5130);
	dataBufferOut(6031) <= dataBufferIn(2057) when (flag_long='1') else dataBufferIn(5213);
	dataBufferOut(6032) <= dataBufferIn(2800) when (flag_long='1') else dataBufferIn(5296);
	dataBufferOut(6033) <= dataBufferIn(3543) when (flag_long='1') else dataBufferIn(5379);
	dataBufferOut(6034) <= dataBufferIn(4286) when (flag_long='1') else dataBufferIn(5462);
	dataBufferOut(6035) <= dataBufferIn(5029) when (flag_long='1') else dataBufferIn(5545);
	dataBufferOut(6036) <= dataBufferIn(5772) when (flag_long='1') else dataBufferIn(5628);
	dataBufferOut(6037) <= dataBufferIn( 371) when (flag_long='1') else dataBufferIn(5711);
	dataBufferOut(6038) <= dataBufferIn(1114) when (flag_long='1') else dataBufferIn(5794);
	dataBufferOut(6039) <= dataBufferIn(1857) when (flag_long='1') else dataBufferIn(5877);
	dataBufferOut(6040) <= dataBufferIn(2600) when (flag_long='1') else dataBufferIn(5960);
	dataBufferOut(6041) <= dataBufferIn(3343) when (flag_long='1') else dataBufferIn(6043);
	dataBufferOut(6042) <= dataBufferIn(4086) when (flag_long='1') else dataBufferIn(6126);
	dataBufferOut(6043) <= dataBufferIn(4829) when (flag_long='1') else dataBufferIn(5153);
	dataBufferOut(6044) <= dataBufferIn(5572) when (flag_long='1') else dataBufferIn(5236);
	dataBufferOut(6045) <= dataBufferIn( 171) when (flag_long='1') else dataBufferIn(5319);
	dataBufferOut(6046) <= dataBufferIn( 914) when (flag_long='1') else dataBufferIn(5402);
	dataBufferOut(6047) <= dataBufferIn(1657) when (flag_long='1') else dataBufferIn(5485);
	dataBufferOut(6048) <= dataBufferIn(2400) when (flag_long='1') else dataBufferIn(5568);
	dataBufferOut(6049) <= dataBufferIn(3143) when (flag_long='1') else dataBufferIn(5651);
	dataBufferOut(6050) <= dataBufferIn(3886) when (flag_long='1') else dataBufferIn(5734);
	dataBufferOut(6051) <= dataBufferIn(4629) when (flag_long='1') else dataBufferIn(5817);
	dataBufferOut(6052) <= dataBufferIn(5372) when (flag_long='1') else dataBufferIn(5900);
	dataBufferOut(6053) <= dataBufferIn(6115) when (flag_long='1') else dataBufferIn(5983);
	dataBufferOut(6054) <= dataBufferIn( 714) when (flag_long='1') else dataBufferIn(6066);
	dataBufferOut(6055) <= dataBufferIn(1457) when (flag_long='1') else dataBufferIn(5093);
	dataBufferOut(6056) <= dataBufferIn(2200) when (flag_long='1') else dataBufferIn(5176);
	dataBufferOut(6057) <= dataBufferIn(2943) when (flag_long='1') else dataBufferIn(5259);
	dataBufferOut(6058) <= dataBufferIn(3686) when (flag_long='1') else dataBufferIn(5342);
	dataBufferOut(6059) <= dataBufferIn(4429) when (flag_long='1') else dataBufferIn(5425);
	dataBufferOut(6060) <= dataBufferIn(5172) when (flag_long='1') else dataBufferIn(5508);
	dataBufferOut(6061) <= dataBufferIn(5915) when (flag_long='1') else dataBufferIn(5591);
	dataBufferOut(6062) <= dataBufferIn( 514) when (flag_long='1') else dataBufferIn(5674);
	dataBufferOut(6063) <= dataBufferIn(1257) when (flag_long='1') else dataBufferIn(5757);
	dataBufferOut(6064) <= dataBufferIn(2000) when (flag_long='1') else dataBufferIn(5840);
	dataBufferOut(6065) <= dataBufferIn(2743) when (flag_long='1') else dataBufferIn(5923);
	dataBufferOut(6066) <= dataBufferIn(3486) when (flag_long='1') else dataBufferIn(6006);
	dataBufferOut(6067) <= dataBufferIn(4229) when (flag_long='1') else dataBufferIn(6089);
	dataBufferOut(6068) <= dataBufferIn(4972) when (flag_long='1') else dataBufferIn(5116);
	dataBufferOut(6069) <= dataBufferIn(5715) when (flag_long='1') else dataBufferIn(5199);
	dataBufferOut(6070) <= dataBufferIn( 314) when (flag_long='1') else dataBufferIn(5282);
	dataBufferOut(6071) <= dataBufferIn(1057) when (flag_long='1') else dataBufferIn(5365);
	dataBufferOut(6072) <= dataBufferIn(1800) when (flag_long='1') else dataBufferIn(5448);
	dataBufferOut(6073) <= dataBufferIn(2543) when (flag_long='1') else dataBufferIn(5531);
	dataBufferOut(6074) <= dataBufferIn(3286) when (flag_long='1') else dataBufferIn(5614);
	dataBufferOut(6075) <= dataBufferIn(4029) when (flag_long='1') else dataBufferIn(5697);
	dataBufferOut(6076) <= dataBufferIn(4772) when (flag_long='1') else dataBufferIn(5780);
	dataBufferOut(6077) <= dataBufferIn(5515) when (flag_long='1') else dataBufferIn(5863);
	dataBufferOut(6078) <= dataBufferIn( 114) when (flag_long='1') else dataBufferIn(5946);
	dataBufferOut(6079) <= dataBufferIn( 857) when (flag_long='1') else dataBufferIn(6029);
	dataBufferOut(6080) <= dataBufferIn(1600) when (flag_long='1') else dataBufferIn(6112);
	dataBufferOut(6081) <= dataBufferIn(2343) when (flag_long='1') else dataBufferIn(5139);
	dataBufferOut(6082) <= dataBufferIn(3086) when (flag_long='1') else dataBufferIn(5222);
	dataBufferOut(6083) <= dataBufferIn(3829) when (flag_long='1') else dataBufferIn(5305);
	dataBufferOut(6084) <= dataBufferIn(4572) when (flag_long='1') else dataBufferIn(5388);
	dataBufferOut(6085) <= dataBufferIn(5315) when (flag_long='1') else dataBufferIn(5471);
	dataBufferOut(6086) <= dataBufferIn(6058) when (flag_long='1') else dataBufferIn(5554);
	dataBufferOut(6087) <= dataBufferIn( 657) when (flag_long='1') else dataBufferIn(5637);
	dataBufferOut(6088) <= dataBufferIn(1400) when (flag_long='1') else dataBufferIn(5720);
	dataBufferOut(6089) <= dataBufferIn(2143) when (flag_long='1') else dataBufferIn(5803);
	dataBufferOut(6090) <= dataBufferIn(2886) when (flag_long='1') else dataBufferIn(5886);
	dataBufferOut(6091) <= dataBufferIn(3629) when (flag_long='1') else dataBufferIn(5969);
	dataBufferOut(6092) <= dataBufferIn(4372) when (flag_long='1') else dataBufferIn(6052);
	dataBufferOut(6093) <= dataBufferIn(5115) when (flag_long='1') else dataBufferIn(6135);
	dataBufferOut(6094) <= dataBufferIn(5858) when (flag_long='1') else dataBufferIn(5162);
	dataBufferOut(6095) <= dataBufferIn( 457) when (flag_long='1') else dataBufferIn(5245);
	dataBufferOut(6096) <= dataBufferIn(1200) when (flag_long='1') else dataBufferIn(5328);
	dataBufferOut(6097) <= dataBufferIn(1943) when (flag_long='1') else dataBufferIn(5411);
	dataBufferOut(6098) <= dataBufferIn(2686) when (flag_long='1') else dataBufferIn(5494);
	dataBufferOut(6099) <= dataBufferIn(3429) when (flag_long='1') else dataBufferIn(5577);
	dataBufferOut(6100) <= dataBufferIn(4172) when (flag_long='1') else dataBufferIn(5660);
	dataBufferOut(6101) <= dataBufferIn(4915) when (flag_long='1') else dataBufferIn(5743);
	dataBufferOut(6102) <= dataBufferIn(5658) when (flag_long='1') else dataBufferIn(5826);
	dataBufferOut(6103) <= dataBufferIn( 257) when (flag_long='1') else dataBufferIn(5909);
	dataBufferOut(6104) <= dataBufferIn(1000) when (flag_long='1') else dataBufferIn(5992);
	dataBufferOut(6105) <= dataBufferIn(1743) when (flag_long='1') else dataBufferIn(6075);
	dataBufferOut(6106) <= dataBufferIn(2486) when (flag_long='1') else dataBufferIn(5102);
	dataBufferOut(6107) <= dataBufferIn(3229) when (flag_long='1') else dataBufferIn(5185);
	dataBufferOut(6108) <= dataBufferIn(3972) when (flag_long='1') else dataBufferIn(5268);
	dataBufferOut(6109) <= dataBufferIn(4715) when (flag_long='1') else dataBufferIn(5351);
	dataBufferOut(6110) <= dataBufferIn(5458) when (flag_long='1') else dataBufferIn(5434);
	dataBufferOut(6111) <= dataBufferIn(  57) when (flag_long='1') else dataBufferIn(5517);
	dataBufferOut(6112) <= dataBufferIn( 800) when (flag_long='1') else dataBufferIn(5600);
	dataBufferOut(6113) <= dataBufferIn(1543) when (flag_long='1') else dataBufferIn(5683);
	dataBufferOut(6114) <= dataBufferIn(2286) when (flag_long='1') else dataBufferIn(5766);
	dataBufferOut(6115) <= dataBufferIn(3029) when (flag_long='1') else dataBufferIn(5849);
	dataBufferOut(6116) <= dataBufferIn(3772) when (flag_long='1') else dataBufferIn(5932);
	dataBufferOut(6117) <= dataBufferIn(4515) when (flag_long='1') else dataBufferIn(6015);
	dataBufferOut(6118) <= dataBufferIn(5258) when (flag_long='1') else dataBufferIn(6098);
	dataBufferOut(6119) <= dataBufferIn(6001) when (flag_long='1') else dataBufferIn(5125);
	dataBufferOut(6120) <= dataBufferIn( 600) when (flag_long='1') else dataBufferIn(5208);
	dataBufferOut(6121) <= dataBufferIn(1343) when (flag_long='1') else dataBufferIn(5291);
	dataBufferOut(6122) <= dataBufferIn(2086) when (flag_long='1') else dataBufferIn(5374);
	dataBufferOut(6123) <= dataBufferIn(2829) when (flag_long='1') else dataBufferIn(5457);
	dataBufferOut(6124) <= dataBufferIn(3572) when (flag_long='1') else dataBufferIn(5540);
	dataBufferOut(6125) <= dataBufferIn(4315) when (flag_long='1') else dataBufferIn(5623);
	dataBufferOut(6126) <= dataBufferIn(5058) when (flag_long='1') else dataBufferIn(5706);
	dataBufferOut(6127) <= dataBufferIn(5801) when (flag_long='1') else dataBufferIn(5789);
	dataBufferOut(6128) <= dataBufferIn( 400) when (flag_long='1') else dataBufferIn(5872);
	dataBufferOut(6129) <= dataBufferIn(1143) when (flag_long='1') else dataBufferIn(5955);
	dataBufferOut(6130) <= dataBufferIn(1886) when (flag_long='1') else dataBufferIn(6038);
	dataBufferOut(6131) <= dataBufferIn(2629) when (flag_long='1') else dataBufferIn(6121);
	dataBufferOut(6132) <= dataBufferIn(3372) when (flag_long='1') else dataBufferIn(5148);
	dataBufferOut(6133) <= dataBufferIn(4115) when (flag_long='1') else dataBufferIn(5231);
	dataBufferOut(6134) <= dataBufferIn(4858) when (flag_long='1') else dataBufferIn(5314);
	dataBufferOut(6135) <= dataBufferIn(5601) when (flag_long='1') else dataBufferIn(5397);
	dataBufferOut(6136) <= dataBufferIn( 200) when (flag_long='1') else dataBufferIn(5480);
	dataBufferOut(6137) <= dataBufferIn( 943) when (flag_long='1') else dataBufferIn(5563);
	dataBufferOut(6138) <= dataBufferIn(1686) when (flag_long='1') else dataBufferIn(5646);
	dataBufferOut(6139) <= dataBufferIn(2429) when (flag_long='1') else dataBufferIn(5729);
	dataBufferOut(6140) <= dataBufferIn(3172) when (flag_long='1') else dataBufferIn(5812);
	dataBufferOut(6141) <= dataBufferIn(3915) when (flag_long='1') else dataBufferIn(5895);
	dataBufferOut(6142) <= dataBufferIn(4658) when (flag_long='1') else dataBufferIn(5978);
	dataBufferOut(6143) <= dataBufferIn(5401) when (flag_long='1') else dataBufferIn(6061);


end arch1;

delay1_inst : delay1 PORT MAP (
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		shiftout	 => shiftout_sig
	);
